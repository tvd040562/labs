module cust_rom1 (clk0,
    cs0,
    addr0,
    dout0);
 input clk0;
 input cs0;
 input [7:0] addr0;
 output [31:0] dout0;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire \addr0_reg[0] ;
 wire \addr0_reg[1] ;
 wire \addr0_reg[2] ;
 wire \addr0_reg[3] ;
 wire \addr0_reg[4] ;
 wire \addr0_reg[5] ;
 wire \addr0_reg[6] ;
 wire \addr0_reg[7] ;
 wire cs0_reg;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire clknet_0_clk0;
 wire clknet_2_0__leaf_clk0;
 wire clknet_2_1__leaf_clk0;
 wire clknet_2_2__leaf_clk0;
 wire clknet_2_3__leaf_clk0;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;

 sky130_fd_sc_hd__inv_2 _0691_ (.A(cs0_reg),
    .Y(_0628_));
 sky130_fd_sc_hd__and4b_1 _0692_ (.A_N(net584),
    .B(net594),
    .C(net600),
    .D(net607),
    .X(_0638_));
 sky130_fd_sc_hd__and4bb_1 _0693_ (.A_N(net558),
    .B_N(net564),
    .C(net570),
    .D(net577),
    .X(_0648_));
 sky130_fd_sc_hd__and4bb_1 _0694_ (.A_N(net600),
    .B_N(net593),
    .C(net584),
    .D(net608),
    .X(_0658_));
 sky130_fd_sc_hd__and4bb_1 _0695_ (.A_N(net570),
    .B_N(net577),
    .C(net558),
    .D(net564),
    .X(_0666_));
 sky130_fd_sc_hd__a22o_1 _0696_ (.A1(net538),
    .A2(net531),
    .B1(net526),
    .B2(net518),
    .X(_0668_));
 sky130_fd_sc_hd__and4bb_1 _0697_ (.A_N(net607),
    .B_N(net585),
    .C(net595),
    .D(net601),
    .X(_0669_));
 sky130_fd_sc_hd__and4bb_1 _0698_ (.A_N(net607),
    .B_N(net593),
    .C(net587),
    .D(net601),
    .X(_0670_));
 sky130_fd_sc_hd__a22o_1 _0699_ (.A1(net530),
    .A2(net514),
    .B1(net507),
    .B2(net519),
    .X(_0671_));
 sky130_fd_sc_hd__and4bb_1 _0700_ (.A_N(net600),
    .B_N(net584),
    .C(net595),
    .D(net610),
    .X(_0672_));
 sky130_fd_sc_hd__and4b_1 _0701_ (.A_N(net593),
    .B(net585),
    .C(net608),
    .D(net601),
    .X(_0673_));
 sky130_fd_sc_hd__a22o_1 _0702_ (.A1(net530),
    .A2(net498),
    .B1(net495),
    .B2(net519),
    .X(_0674_));
 sky130_fd_sc_hd__or4b_1 _0703_ (.A(net600),
    .B(net607),
    .C(net593),
    .D_N(net584),
    .X(_0675_));
 sky130_fd_sc_hd__o21ba_1 _0704_ (.A1(net530),
    .A2(net518),
    .B1_N(net489),
    .X(_0676_));
 sky130_fd_sc_hd__or3_1 _0705_ (.A(net331),
    .B(net327),
    .C(net324),
    .X(_0677_));
 sky130_fd_sc_hd__or4_1 _0706_ (.A(net334),
    .B(net332),
    .C(net327),
    .D(net324),
    .X(_0678_));
 sky130_fd_sc_hd__and4b_1 _0707_ (.A_N(net612),
    .B(net590),
    .C(net599),
    .D(net603),
    .X(_0679_));
 sky130_fd_sc_hd__nor4b_1 _0708_ (.A(net612),
    .B(net589),
    .C(net597),
    .D_N(net604),
    .Y(_0680_));
 sky130_fd_sc_hd__a22o_1 _0709_ (.A1(net532),
    .A2(net482),
    .B1(net475),
    .B2(net520),
    .X(_0681_));
 sky130_fd_sc_hd__and4_1 _0710_ (.A(net603),
    .B(net612),
    .C(net589),
    .D(net597),
    .X(_0682_));
 sky130_fd_sc_hd__nor4b_1 _0711_ (.A(net603),
    .B(net589),
    .C(net597),
    .D_N(net612),
    .Y(_0683_));
 sky130_fd_sc_hd__a22o_1 _0712_ (.A1(net532),
    .A2(net467),
    .B1(net459),
    .B2(net520),
    .X(_0684_));
 sky130_fd_sc_hd__or2_1 _0713_ (.A(net323),
    .B(net318),
    .X(_0685_));
 sky130_fd_sc_hd__or4_1 _0714_ (.A(net605),
    .B(net614),
    .C(net591),
    .D(net598),
    .X(_0686_));
 sky130_fd_sc_hd__nor4b_1 _0715_ (.A(net575),
    .B(net457),
    .C(net582),
    .D_N(net568),
    .Y(_0687_));
 sky130_fd_sc_hd__and4b_1 _0716_ (.A_N(net602),
    .B(net611),
    .C(net588),
    .D(net596),
    .X(_0688_));
 sky130_fd_sc_hd__and4bb_1 _0717_ (.A_N(net589),
    .B_N(net597),
    .C(net603),
    .D(net613),
    .X(_0689_));
 sky130_fd_sc_hd__a22o_1 _0718_ (.A1(net531),
    .A2(net450),
    .B1(net443),
    .B2(net518),
    .X(_0690_));
 sky130_fd_sc_hd__or2_1 _0719_ (.A(net322),
    .B(net315),
    .X(_0031_));
 sky130_fd_sc_hd__or3_1 _0720_ (.A(net323),
    .B(net318),
    .C(net316),
    .X(_0032_));
 sky130_fd_sc_hd__or4_1 _0721_ (.A(net322),
    .B(net318),
    .C(net316),
    .D(net314),
    .X(_0033_));
 sky130_fd_sc_hd__and4bb_1 _0722_ (.A_N(net605),
    .B_N(net614),
    .C(net591),
    .D(net598),
    .X(_0034_));
 sky130_fd_sc_hd__nor4b_1 _0723_ (.A(net605),
    .B(net614),
    .C(net591),
    .D_N(net598),
    .Y(_0035_));
 sky130_fd_sc_hd__a22o_1 _0724_ (.A1(net534),
    .A2(net438),
    .B1(net431),
    .B2(net519),
    .X(_0036_));
 sky130_fd_sc_hd__a22o_1 _0725_ (.A1(net531),
    .A2(net526),
    .B1(net518),
    .B2(net538),
    .X(_0037_));
 sky130_fd_sc_hd__a22o_1 _0726_ (.A1(net521),
    .A2(net511),
    .B1(net504),
    .B2(net533),
    .X(_0038_));
 sky130_fd_sc_hd__a22o_1 _0727_ (.A1(net521),
    .A2(net499),
    .B1(net491),
    .B2(net533),
    .X(_0039_));
 sky130_fd_sc_hd__or3_2 _0728_ (.A(_0037_),
    .B(net309),
    .C(net308),
    .X(_0040_));
 sky130_fd_sc_hd__or2_1 _0729_ (.A(net312),
    .B(net307),
    .X(_0041_));
 sky130_fd_sc_hd__or4_1 _0730_ (.A(net312),
    .B(net310),
    .C(net309),
    .D(net307),
    .X(_0042_));
 sky130_fd_sc_hd__a22o_1 _0731_ (.A1(net521),
    .A2(net450),
    .B1(net443),
    .B2(net533),
    .X(_0043_));
 sky130_fd_sc_hd__a22o_1 _0732_ (.A1(net520),
    .A2(net436),
    .B1(net430),
    .B2(net532),
    .X(_0044_));
 sky130_fd_sc_hd__a22o_1 _0733_ (.A1(net520),
    .A2(net467),
    .B1(net459),
    .B2(net532),
    .X(_0045_));
 sky130_fd_sc_hd__a22o_1 _0734_ (.A1(net521),
    .A2(net483),
    .B1(net476),
    .B2(net533),
    .X(_0046_));
 sky130_fd_sc_hd__or2_1 _0735_ (.A(net304),
    .B(net298),
    .X(_0047_));
 sky130_fd_sc_hd__or3_1 _0736_ (.A(net304),
    .B(net301),
    .C(net296),
    .X(_0048_));
 sky130_fd_sc_hd__or2_1 _0737_ (.A(net305),
    .B(net300),
    .X(_0049_));
 sky130_fd_sc_hd__or4_1 _0738_ (.A(net305),
    .B(_0044_),
    .C(net300),
    .D(net297),
    .X(_0050_));
 sky130_fd_sc_hd__or4_1 _0739_ (.A(_0678_),
    .B(_0033_),
    .C(_0042_),
    .D(_0050_),
    .X(_0051_));
 sky130_fd_sc_hd__and4bb_1 _0740_ (.A_N(net579),
    .B_N(net559),
    .C(net565),
    .D(net572),
    .X(_0052_));
 sky130_fd_sc_hd__and4bb_1 _0741_ (.A_N(net570),
    .B_N(net564),
    .C(net558),
    .D(net577),
    .X(_0053_));
 sky130_fd_sc_hd__a22o_1 _0742_ (.A1(net535),
    .A2(net422),
    .B1(net415),
    .B2(net523),
    .X(_0054_));
 sky130_fd_sc_hd__a22o_1 _0743_ (.A1(net499),
    .A2(net422),
    .B1(net415),
    .B2(net492),
    .X(_0055_));
 sky130_fd_sc_hd__o21ba_1 _0744_ (.A1(net422),
    .A2(net415),
    .B1_N(net490),
    .X(_0056_));
 sky130_fd_sc_hd__a22o_1 _0745_ (.A1(net512),
    .A2(net424),
    .B1(net417),
    .B2(net505),
    .X(_0057_));
 sky130_fd_sc_hd__or2_1 _0746_ (.A(net291),
    .B(net289),
    .X(_0058_));
 sky130_fd_sc_hd__or2_1 _0747_ (.A(net293),
    .B(net289),
    .X(_0059_));
 sky130_fd_sc_hd__or3_2 _0748_ (.A(net295),
    .B(net292),
    .C(net288),
    .X(_0060_));
 sky130_fd_sc_hd__or4_1 _0749_ (.A(net295),
    .B(net292),
    .C(net290),
    .D(net288),
    .X(_0061_));
 sky130_fd_sc_hd__a22o_1 _0750_ (.A1(net491),
    .A2(net423),
    .B1(net416),
    .B2(net499),
    .X(_0062_));
 sky130_fd_sc_hd__a22o_1 _0751_ (.A1(net509),
    .A2(net426),
    .B1(net420),
    .B2(net516),
    .X(_0063_));
 sky130_fd_sc_hd__or2_1 _0752_ (.A(net287),
    .B(net285),
    .X(_0064_));
 sky130_fd_sc_hd__a22o_1 _0753_ (.A1(net524),
    .A2(net422),
    .B1(net415),
    .B2(net536),
    .X(_0065_));
 sky130_fd_sc_hd__or3_1 _0754_ (.A(_0061_),
    .B(_0064_),
    .C(net282),
    .X(_0066_));
 sky130_fd_sc_hd__and4bb_1 _0755_ (.A_N(net574),
    .B_N(net561),
    .C(net567),
    .D(net581),
    .X(_0067_));
 sky130_fd_sc_hd__and4bb_1 _0756_ (.A_N(net581),
    .B_N(net567),
    .C(net561),
    .D(net574),
    .X(_0068_));
 sky130_fd_sc_hd__a22o_1 _0757_ (.A1(net496),
    .A2(net409),
    .B1(net400),
    .B2(net503),
    .X(_0069_));
 sky130_fd_sc_hd__a22o_1 _0758_ (.A1(net441),
    .A2(net412),
    .B1(net403),
    .B2(net434),
    .X(_0070_));
 sky130_fd_sc_hd__a22o_1 _0759_ (.A1(net527),
    .A2(net409),
    .B1(net400),
    .B2(net539),
    .X(_0071_));
 sky130_fd_sc_hd__a22o_1 _0760_ (.A1(net509),
    .A2(net411),
    .B1(net402),
    .B2(net516),
    .X(_0072_));
 sky130_fd_sc_hd__or2_1 _0761_ (.A(_0071_),
    .B(net277),
    .X(_0073_));
 sky130_fd_sc_hd__or3_2 _0762_ (.A(net281),
    .B(net279),
    .C(net276),
    .X(_0074_));
 sky130_fd_sc_hd__or4_2 _0763_ (.A(net280),
    .B(_0070_),
    .C(net278),
    .D(net276),
    .X(_0075_));
 sky130_fd_sc_hd__a22o_1 _0764_ (.A1(net484),
    .A2(net408),
    .B1(net399),
    .B2(net477),
    .X(_0076_));
 sky130_fd_sc_hd__a22o_1 _0765_ (.A1(net453),
    .A2(net406),
    .B1(net398),
    .B2(net446),
    .X(_0077_));
 sky130_fd_sc_hd__a22o_1 _0766_ (.A1(net473),
    .A2(net410),
    .B1(net401),
    .B2(net465),
    .X(_0078_));
 sky130_fd_sc_hd__o21ba_1 _0767_ (.A1(net426),
    .A2(net402),
    .B1_N(net458),
    .X(_0079_));
 sky130_fd_sc_hd__or2_1 _0768_ (.A(net270),
    .B(net269),
    .X(_0080_));
 sky130_fd_sc_hd__or4_1 _0769_ (.A(_0075_),
    .B(net272),
    .C(net271),
    .D(_0080_),
    .X(_0081_));
 sky130_fd_sc_hd__and4b_1 _0770_ (.A_N(net561),
    .B(net567),
    .C(net574),
    .D(net581),
    .X(_0082_));
 sky130_fd_sc_hd__nor4b_1 _0771_ (.A(net575),
    .B(net581),
    .C(net567),
    .D_N(net561),
    .Y(_0083_));
 sky130_fd_sc_hd__a22o_1 _0772_ (.A1(net446),
    .A2(net392),
    .B1(net386),
    .B2(net453),
    .X(_0084_));
 sky130_fd_sc_hd__a22o_1 _0773_ (.A1(net433),
    .A2(net393),
    .B1(net387),
    .B2(net440),
    .X(_0085_));
 sky130_fd_sc_hd__a22o_1 _0774_ (.A1(net461),
    .A2(net392),
    .B1(net386),
    .B2(net469),
    .X(_0086_));
 sky130_fd_sc_hd__a22o_1 _0775_ (.A1(net477),
    .A2(net392),
    .B1(net386),
    .B2(net484),
    .X(_0087_));
 sky130_fd_sc_hd__or2_1 _0776_ (.A(net263),
    .B(net260),
    .X(_0088_));
 sky130_fd_sc_hd__or3_1 _0777_ (.A(net266),
    .B(net264),
    .C(net260),
    .X(_0089_));
 sky130_fd_sc_hd__or4_1 _0778_ (.A(net266),
    .B(net264),
    .C(net263),
    .D(net260),
    .X(_0090_));
 sky130_fd_sc_hd__a22o_1 _0779_ (.A1(_0672_),
    .A2(net394),
    .B1(net388),
    .B2(net497),
    .X(_0091_));
 sky130_fd_sc_hd__a22o_1 _0780_ (.A1(net539),
    .A2(net396),
    .B1(net390),
    .B2(net527),
    .X(_0092_));
 sky130_fd_sc_hd__or2_1 _0781_ (.A(net258),
    .B(net256),
    .X(_0093_));
 sky130_fd_sc_hd__o21ba_1 _0782_ (.A1(net392),
    .A2(net386),
    .B1_N(net489),
    .X(_0094_));
 sky130_fd_sc_hd__a22o_1 _0783_ (.A1(net515),
    .A2(net396),
    .B1(net390),
    .B2(net508),
    .X(_0095_));
 sky130_fd_sc_hd__or2_1 _0784_ (.A(net254),
    .B(net253),
    .X(_0096_));
 sky130_fd_sc_hd__or4_1 _0785_ (.A(net258),
    .B(net256),
    .C(net254),
    .D(net252),
    .X(_0097_));
 sky130_fd_sc_hd__or2_1 _0786_ (.A(_0090_),
    .B(_0097_),
    .X(_0098_));
 sky130_fd_sc_hd__nor4b_1 _0787_ (.A(net570),
    .B(net577),
    .C(net558),
    .D_N(net565),
    .Y(_0099_));
 sky130_fd_sc_hd__and4b_1 _0788_ (.A_N(net566),
    .B(net560),
    .C(net580),
    .D(net573),
    .X(_0100_));
 sky130_fd_sc_hd__o21ba_1 _0789_ (.A1(net380),
    .A2(net374),
    .B1_N(net490),
    .X(_0101_));
 sky130_fd_sc_hd__a22o_1 _0790_ (.A1(net535),
    .A2(net380),
    .B1(net374),
    .B2(net523),
    .X(_0102_));
 sky130_fd_sc_hd__or2_1 _0791_ (.A(net250),
    .B(net249),
    .X(_0103_));
 sky130_fd_sc_hd__a22o_1 _0792_ (.A1(net500),
    .A2(net384),
    .B1(net376),
    .B2(net491),
    .X(_0104_));
 sky130_fd_sc_hd__a22o_1 _0793_ (.A1(net512),
    .A2(net382),
    .B1(net376),
    .B2(net504),
    .X(_0105_));
 sky130_fd_sc_hd__or2_1 _0794_ (.A(net247),
    .B(net245),
    .X(_0106_));
 sky130_fd_sc_hd__or4_2 _0795_ (.A(net250),
    .B(net248),
    .C(net246),
    .D(net245),
    .X(_0107_));
 sky130_fd_sc_hd__o21ba_1 _0796_ (.A1(net413),
    .A2(net404),
    .B1_N(net489),
    .X(_0108_));
 sky130_fd_sc_hd__a22o_1 _0797_ (.A1(net539),
    .A2(net409),
    .B1(net400),
    .B2(net527),
    .X(_0109_));
 sky130_fd_sc_hd__or2_1 _0798_ (.A(net242),
    .B(net241),
    .X(_0110_));
 sky130_fd_sc_hd__a22o_1 _0799_ (.A1(net513),
    .A2(net406),
    .B1(net398),
    .B2(net506),
    .X(_0111_));
 sky130_fd_sc_hd__a22o_1 _0800_ (.A1(net503),
    .A2(net406),
    .B1(net398),
    .B2(net496),
    .X(_0112_));
 sky130_fd_sc_hd__or2_1 _0801_ (.A(net238),
    .B(_0112_),
    .X(_0113_));
 sky130_fd_sc_hd__or2_2 _0802_ (.A(net240),
    .B(_0112_),
    .X(_0114_));
 sky130_fd_sc_hd__or3_1 _0803_ (.A(_0107_),
    .B(net63),
    .C(_0113_),
    .X(_0115_));
 sky130_fd_sc_hd__nor4b_1 _0804_ (.A(net580),
    .B(net560),
    .C(net566),
    .D_N(net573),
    .Y(_0116_));
 sky130_fd_sc_hd__and4b_1 _0805_ (.A_N(net571),
    .B(net578),
    .C(net559),
    .D(net564),
    .X(_0117_));
 sky130_fd_sc_hd__a22o_1 _0806_ (.A1(net476),
    .A2(net367),
    .B1(net361),
    .B2(net483),
    .X(_0118_));
 sky130_fd_sc_hd__a22o_1 _0807_ (.A1(net459),
    .A2(net371),
    .B1(net365),
    .B2(net467),
    .X(_0119_));
 sky130_fd_sc_hd__a22o_1 _0808_ (.A1(net444),
    .A2(net367),
    .B1(net361),
    .B2(net451),
    .X(_0120_));
 sky130_fd_sc_hd__a22o_1 _0809_ (.A1(net429),
    .A2(net367),
    .B1(net361),
    .B2(net437),
    .X(_0121_));
 sky130_fd_sc_hd__or2_1 _0810_ (.A(net232),
    .B(net228),
    .X(_0122_));
 sky130_fd_sc_hd__or4_2 _0811_ (.A(net236),
    .B(net235),
    .C(net231),
    .D(net230),
    .X(_0123_));
 sky130_fd_sc_hd__a22o_1 _0812_ (.A1(net511),
    .A2(net369),
    .B1(net363),
    .B2(net505),
    .X(_0124_));
 sky130_fd_sc_hd__a22o_1 _0813_ (.A1(net499),
    .A2(net369),
    .B1(net363),
    .B2(net491),
    .X(_0125_));
 sky130_fd_sc_hd__o21ba_1 _0814_ (.A1(net370),
    .A2(net364),
    .B1_N(net490),
    .X(_0126_));
 sky130_fd_sc_hd__a22o_1 _0815_ (.A1(net537),
    .A2(net370),
    .B1(net364),
    .B2(net525),
    .X(_0127_));
 sky130_fd_sc_hd__or3_1 _0816_ (.A(net225),
    .B(net224),
    .C(net218),
    .X(_0128_));
 sky130_fd_sc_hd__or4_1 _0817_ (.A(net226),
    .B(net224),
    .C(net221),
    .D(net219),
    .X(_0129_));
 sky130_fd_sc_hd__or2_1 _0818_ (.A(net62),
    .B(_0129_),
    .X(_0130_));
 sky130_fd_sc_hd__a22o_1 _0819_ (.A1(net495),
    .A2(net368),
    .B1(net362),
    .B2(net498),
    .X(_0131_));
 sky130_fd_sc_hd__a22o_1 _0820_ (.A1(net437),
    .A2(net367),
    .B1(net361),
    .B2(net429),
    .X(_0132_));
 sky130_fd_sc_hd__a22o_1 _0821_ (.A1(net497),
    .A2(net394),
    .B1(net388),
    .B2(net503),
    .X(_0133_));
 sky130_fd_sc_hd__a22o_1 _0822_ (.A1(net440),
    .A2(net395),
    .B1(net387),
    .B2(net433),
    .X(_0134_));
 sky130_fd_sc_hd__or2_1 _0823_ (.A(_0133_),
    .B(net210),
    .X(_0135_));
 sky130_fd_sc_hd__and2b_1 _0824_ (.A_N(net458),
    .B(net389),
    .X(_0136_));
 sky130_fd_sc_hd__a22o_1 _0825_ (.A1(net439),
    .A2(net426),
    .B1(net420),
    .B2(net432),
    .X(_0137_));
 sky130_fd_sc_hd__a22o_1 _0826_ (.A1(net527),
    .A2(net394),
    .B1(net388),
    .B2(net539),
    .X(_0138_));
 sky130_fd_sc_hd__a22o_1 _0827_ (.A1(net509),
    .A2(net396),
    .B1(net390),
    .B2(net516),
    .X(_0139_));
 sky130_fd_sc_hd__a22o_1 _0828_ (.A1(net523),
    .A2(net371),
    .B1(net365),
    .B2(net535),
    .X(_0140_));
 sky130_fd_sc_hd__a22o_1 _0829_ (.A1(net504),
    .A2(net369),
    .B1(net363),
    .B2(net511),
    .X(_0141_));
 sky130_fd_sc_hd__or4_1 _0830_ (.A(net206),
    .B(net205),
    .C(net202),
    .D(net199),
    .X(_0142_));
 sky130_fd_sc_hd__o21ba_1 _0831_ (.A1(net419),
    .A2(net393),
    .B1_N(net458),
    .X(_0143_));
 sky130_fd_sc_hd__a22o_1 _0832_ (.A1(net483),
    .A2(net425),
    .B1(net418),
    .B2(net476),
    .X(_0144_));
 sky130_fd_sc_hd__a22o_1 _0833_ (.A1(net451),
    .A2(net423),
    .B1(net416),
    .B2(net444),
    .X(_0145_));
 sky130_fd_sc_hd__a22o_1 _0834_ (.A1(net470),
    .A2(net427),
    .B1(net420),
    .B2(net462),
    .X(_0146_));
 sky130_fd_sc_hd__or2_1 _0835_ (.A(net194),
    .B(net191),
    .X(_0147_));
 sky130_fd_sc_hd__or2_1 _0836_ (.A(net198),
    .B(net194),
    .X(_0148_));
 sky130_fd_sc_hd__or4_1 _0837_ (.A(net197),
    .B(net196),
    .C(net193),
    .D(net191),
    .X(_0149_));
 sky130_fd_sc_hd__nor4_1 _0838_ (.A(net575),
    .B(net582),
    .C(net562),
    .D(net568),
    .Y(_0150_));
 sky130_fd_sc_hd__and4_1 _0839_ (.A(net574),
    .B(net582),
    .C(net562),
    .D(net568),
    .X(_0151_));
 sky130_fd_sc_hd__a22o_1 _0840_ (.A1(net432),
    .A2(net359),
    .B1(net349),
    .B2(net440),
    .X(_0152_));
 sky130_fd_sc_hd__a22o_1 _0841_ (.A1(net478),
    .A2(net357),
    .B1(net351),
    .B2(net485),
    .X(_0153_));
 sky130_fd_sc_hd__a22o_1 _0842_ (.A1(net462),
    .A2(net356),
    .B1(net350),
    .B2(net470),
    .X(_0154_));
 sky130_fd_sc_hd__or2_2 _0843_ (.A(net188),
    .B(net184),
    .X(_0155_));
 sky130_fd_sc_hd__a22o_1 _0844_ (.A1(net448),
    .A2(net356),
    .B1(net350),
    .B2(net454),
    .X(_0156_));
 sky130_fd_sc_hd__or2_1 _0845_ (.A(_0155_),
    .B(net183),
    .X(_0157_));
 sky130_fd_sc_hd__or4_2 _0846_ (.A(net189),
    .B(net187),
    .C(net184),
    .D(net182),
    .X(_0158_));
 sky130_fd_sc_hd__a22o_1 _0847_ (.A1(net515),
    .A2(net355),
    .B1(net348),
    .B2(net508),
    .X(_0159_));
 sky130_fd_sc_hd__o21ba_1 _0848_ (.A1(net360),
    .A2(net354),
    .B1_N(net490),
    .X(_0160_));
 sky130_fd_sc_hd__or2_1 _0849_ (.A(net181),
    .B(net179),
    .X(_0161_));
 sky130_fd_sc_hd__a22o_1 _0850_ (.A1(net498),
    .A2(net360),
    .B1(net354),
    .B2(net495),
    .X(_0162_));
 sky130_fd_sc_hd__a22o_1 _0851_ (.A1(net540),
    .A2(net355),
    .B1(net348),
    .B2(net528),
    .X(_0163_));
 sky130_fd_sc_hd__or4_2 _0852_ (.A(net181),
    .B(net179),
    .C(net177),
    .D(net175),
    .X(_0164_));
 sky130_fd_sc_hd__a22o_1 _0853_ (.A1(net439),
    .A2(net358),
    .B1(net352),
    .B2(net433),
    .X(_0165_));
 sky130_fd_sc_hd__a22o_1 _0854_ (.A1(net494),
    .A2(net360),
    .B1(net354),
    .B2(net502),
    .X(_0166_));
 sky130_fd_sc_hd__a22o_1 _0855_ (.A1(net508),
    .A2(net355),
    .B1(net349),
    .B2(net515),
    .X(_0167_));
 sky130_fd_sc_hd__a22o_1 _0856_ (.A1(net528),
    .A2(net355),
    .B1(net348),
    .B2(net540),
    .X(_0168_));
 sky130_fd_sc_hd__or2_1 _0857_ (.A(_0167_),
    .B(net165),
    .X(_0169_));
 sky130_fd_sc_hd__or2_1 _0858_ (.A(net171),
    .B(net167),
    .X(_0170_));
 sky130_fd_sc_hd__or4_1 _0859_ (.A(net172),
    .B(net169),
    .C(net167),
    .D(net165),
    .X(_0171_));
 sky130_fd_sc_hd__or2_1 _0860_ (.A(_0164_),
    .B(_0171_),
    .X(_0172_));
 sky130_fd_sc_hd__a22o_1 _0861_ (.A1(net470),
    .A2(net356),
    .B1(net350),
    .B2(net462),
    .X(_0173_));
 sky130_fd_sc_hd__a22o_1 _0862_ (.A1(net486),
    .A2(net357),
    .B1(net351),
    .B2(net479),
    .X(_0174_));
 sky130_fd_sc_hd__or2_1 _0863_ (.A(net162),
    .B(net160),
    .X(_0175_));
 sky130_fd_sc_hd__a22o_1 _0864_ (.A1(net455),
    .A2(net356),
    .B1(net350),
    .B2(net447),
    .X(_0176_));
 sky130_fd_sc_hd__nor4b_1 _0865_ (.A(net573),
    .B(net560),
    .C(net566),
    .D_N(net580),
    .Y(_0177_));
 sky130_fd_sc_hd__o21ba_1 _0866_ (.A1(net348),
    .A2(net344),
    .B1_N(net458),
    .X(_0178_));
 sky130_fd_sc_hd__or2_1 _0867_ (.A(net160),
    .B(net157),
    .X(_0179_));
 sky130_fd_sc_hd__or2_1 _0868_ (.A(net162),
    .B(net158),
    .X(_0180_));
 sky130_fd_sc_hd__or2_1 _0869_ (.A(net159),
    .B(net154),
    .X(_0181_));
 sky130_fd_sc_hd__or4_1 _0870_ (.A(net163),
    .B(net159),
    .C(_0176_),
    .D(net154),
    .X(_0182_));
 sky130_fd_sc_hd__or4_1 _0871_ (.A(_0158_),
    .B(_0164_),
    .C(_0171_),
    .D(_0182_),
    .X(_0183_));
 sky130_fd_sc_hd__and4b_1 _0872_ (.A_N(net580),
    .B(net560),
    .C(net566),
    .D(net573),
    .X(_0184_));
 sky130_fd_sc_hd__a22o_1 _0873_ (.A1(net439),
    .A2(net344),
    .B1(net338),
    .B2(net432),
    .X(_0185_));
 sky130_fd_sc_hd__a22o_1 _0874_ (.A1(net507),
    .A2(net342),
    .B1(net335),
    .B2(net514),
    .X(_0186_));
 sky130_fd_sc_hd__a22o_1 _0875_ (.A1(net524),
    .A2(net343),
    .B1(net335),
    .B2(net536),
    .X(_0187_));
 sky130_fd_sc_hd__a22o_1 _0876_ (.A1(net493),
    .A2(net342),
    .B1(net336),
    .B2(net501),
    .X(_0188_));
 sky130_fd_sc_hd__or2_1 _0877_ (.A(net148),
    .B(net147),
    .X(_0189_));
 sky130_fd_sc_hd__or2_1 _0878_ (.A(net151),
    .B(net149),
    .X(_0190_));
 sky130_fd_sc_hd__or3_1 _0879_ (.A(net150),
    .B(net148),
    .C(net146),
    .X(_0191_));
 sky130_fd_sc_hd__or2_2 _0880_ (.A(net152),
    .B(net146),
    .X(_0192_));
 sky130_fd_sc_hd__or2_1 _0881_ (.A(_0190_),
    .B(_0192_),
    .X(_0193_));
 sky130_fd_sc_hd__a22o_1 _0882_ (.A1(net446),
    .A2(net347),
    .B1(net341),
    .B2(net453),
    .X(_0194_));
 sky130_fd_sc_hd__a22o_1 _0883_ (.A1(net432),
    .A2(net344),
    .B1(net339),
    .B2(net439),
    .X(_0195_));
 sky130_fd_sc_hd__a22o_1 _0884_ (.A1(net478),
    .A2(net345),
    .B1(net338),
    .B2(net485),
    .X(_0196_));
 sky130_fd_sc_hd__a22o_1 _0885_ (.A1(net464),
    .A2(net345),
    .B1(net338),
    .B2(net472),
    .X(_0197_));
 sky130_fd_sc_hd__or2_1 _0886_ (.A(net141),
    .B(net140),
    .X(_0198_));
 sky130_fd_sc_hd__or2_1 _0887_ (.A(_0195_),
    .B(net141),
    .X(_0199_));
 sky130_fd_sc_hd__or3_1 _0888_ (.A(net144),
    .B(net141),
    .C(net140),
    .X(_0200_));
 sky130_fd_sc_hd__or4_2 _0889_ (.A(net145),
    .B(net144),
    .C(net141),
    .D(net140),
    .X(_0201_));
 sky130_fd_sc_hd__o21ba_1 _0890_ (.A1(net342),
    .A2(net335),
    .B1_N(net489),
    .X(_0202_));
 sky130_fd_sc_hd__a22o_1 _0891_ (.A1(net515),
    .A2(net343),
    .B1(net337),
    .B2(net508),
    .X(_0203_));
 sky130_fd_sc_hd__or2_2 _0892_ (.A(net137),
    .B(_0203_),
    .X(_0204_));
 sky130_fd_sc_hd__a22o_1 _0893_ (.A1(net538),
    .A2(net342),
    .B1(net335),
    .B2(net526),
    .X(_0205_));
 sky130_fd_sc_hd__a22o_1 _0894_ (.A1(net498),
    .A2(net343),
    .B1(net337),
    .B2(net495),
    .X(_0206_));
 sky130_fd_sc_hd__or2_1 _0895_ (.A(net136),
    .B(net132),
    .X(_0207_));
 sky130_fd_sc_hd__or4_2 _0896_ (.A(net138),
    .B(net136),
    .C(net134),
    .D(net133),
    .X(_0208_));
 sky130_fd_sc_hd__a22o_1 _0897_ (.A1(net486),
    .A2(net344),
    .B1(net339),
    .B2(net479),
    .X(_0209_));
 sky130_fd_sc_hd__a22o_1 _0898_ (.A1(net454),
    .A2(net345),
    .B1(net338),
    .B2(net447),
    .X(_0210_));
 sky130_fd_sc_hd__a22o_1 _0899_ (.A1(net471),
    .A2(net346),
    .B1(net339),
    .B2(net462),
    .X(_0211_));
 sky130_fd_sc_hd__o21ba_1 _0900_ (.A1(net368),
    .A2(net336),
    .B1_N(net457),
    .X(_0212_));
 sky130_fd_sc_hd__or2_1 _0901_ (.A(net127),
    .B(net124),
    .X(_0213_));
 sky130_fd_sc_hd__or2_1 _0902_ (.A(net131),
    .B(net127),
    .X(_0214_));
 sky130_fd_sc_hd__or2_1 _0903_ (.A(net128),
    .B(net124),
    .X(_0215_));
 sky130_fd_sc_hd__or2_1 _0904_ (.A(_0214_),
    .B(_0215_),
    .X(_0216_));
 sky130_fd_sc_hd__or2_1 _0905_ (.A(_0201_),
    .B(_0208_),
    .X(_0217_));
 sky130_fd_sc_hd__or4_1 _0906_ (.A(_0183_),
    .B(_0193_),
    .C(_0216_),
    .D(_0217_),
    .X(_0218_));
 sky130_fd_sc_hd__a22o_1 _0907_ (.A1(net443),
    .A2(net383),
    .B1(net377),
    .B2(net450),
    .X(_0219_));
 sky130_fd_sc_hd__a22o_1 _0908_ (.A1(net459),
    .A2(net379),
    .B1(net373),
    .B2(net467),
    .X(_0220_));
 sky130_fd_sc_hd__or2_1 _0909_ (.A(net123),
    .B(net122),
    .X(_0221_));
 sky130_fd_sc_hd__a22o_1 _0910_ (.A1(net429),
    .A2(net383),
    .B1(net377),
    .B2(net436),
    .X(_0222_));
 sky130_fd_sc_hd__a22o_1 _0911_ (.A1(net475),
    .A2(net379),
    .B1(net373),
    .B2(net482),
    .X(_0223_));
 sky130_fd_sc_hd__or2_1 _0912_ (.A(net119),
    .B(net116),
    .X(_0224_));
 sky130_fd_sc_hd__or4_1 _0913_ (.A(net123),
    .B(_0220_),
    .C(_0222_),
    .D(net117),
    .X(_0225_));
 sky130_fd_sc_hd__a22o_1 _0914_ (.A1(net468),
    .A2(net369),
    .B1(net363),
    .B2(net460),
    .X(_0226_));
 sky130_fd_sc_hd__a22o_1 _0915_ (.A1(net482),
    .A2(net371),
    .B1(net365),
    .B2(net475),
    .X(_0227_));
 sky130_fd_sc_hd__a22o_1 _0916_ (.A1(net450),
    .A2(net368),
    .B1(net362),
    .B2(net443),
    .X(_0228_));
 sky130_fd_sc_hd__o21ba_1 _0917_ (.A1(net530),
    .A2(net362),
    .B1_N(net457),
    .X(_0229_));
 sky130_fd_sc_hd__or3_1 _0918_ (.A(net111),
    .B(net109),
    .C(net104),
    .X(_0230_));
 sky130_fd_sc_hd__or2_1 _0919_ (.A(net113),
    .B(net110),
    .X(_0231_));
 sky130_fd_sc_hd__or4_1 _0920_ (.A(net114),
    .B(net111),
    .C(net109),
    .D(net105),
    .X(_0232_));
 sky130_fd_sc_hd__a22o_1 _0921_ (.A1(net492),
    .A2(net382),
    .B1(net378),
    .B2(net500),
    .X(_0233_));
 sky130_fd_sc_hd__a22o_1 _0922_ (.A1(net523),
    .A2(net379),
    .B1(net373),
    .B2(net535),
    .X(_0234_));
 sky130_fd_sc_hd__a22o_1 _0923_ (.A1(net504),
    .A2(net382),
    .B1(net376),
    .B2(net511),
    .X(_0235_));
 sky130_fd_sc_hd__a22o_1 _0924_ (.A1(net436),
    .A2(net381),
    .B1(net375),
    .B2(net430),
    .X(_0236_));
 sky130_fd_sc_hd__or2_1 _0925_ (.A(net99),
    .B(net96),
    .X(_0237_));
 sky130_fd_sc_hd__or3_1 _0926_ (.A(net102),
    .B(net98),
    .C(net97),
    .X(_0238_));
 sky130_fd_sc_hd__or2_1 _0927_ (.A(net103),
    .B(net96),
    .X(_0239_));
 sky130_fd_sc_hd__or4_1 _0928_ (.A(_0233_),
    .B(net102),
    .C(net99),
    .D(net96),
    .X(_0240_));
 sky130_fd_sc_hd__a22o_1 _0929_ (.A1(net482),
    .A2(net379),
    .B1(net373),
    .B2(net475),
    .X(_0241_));
 sky130_fd_sc_hd__o21ba_1 _0930_ (.A1(net406),
    .A2(net377),
    .B1_N(net457),
    .X(_0242_));
 sky130_fd_sc_hd__or2_2 _0931_ (.A(net95),
    .B(net93),
    .X(_0243_));
 sky130_fd_sc_hd__a22o_1 _0932_ (.A1(net451),
    .A2(net381),
    .B1(net375),
    .B2(net444),
    .X(_0244_));
 sky130_fd_sc_hd__a22o_1 _0933_ (.A1(net468),
    .A2(net383),
    .B1(net377),
    .B2(net460),
    .X(_0245_));
 sky130_fd_sc_hd__or2_2 _0934_ (.A(_0244_),
    .B(net90),
    .X(_0246_));
 sky130_fd_sc_hd__or3_1 _0935_ (.A(_0240_),
    .B(_0243_),
    .C(_0246_),
    .X(_0247_));
 sky130_fd_sc_hd__a22o_1 _0936_ (.A1(net434),
    .A2(net407),
    .B1(net399),
    .B2(net441),
    .X(_0248_));
 sky130_fd_sc_hd__a22o_1 _0937_ (.A1(net448),
    .A2(net409),
    .B1(net400),
    .B2(net455),
    .X(_0249_));
 sky130_fd_sc_hd__or2_1 _0938_ (.A(net89),
    .B(net87),
    .X(_0250_));
 sky130_fd_sc_hd__a22o_1 _0939_ (.A1(net465),
    .A2(net410),
    .B1(net403),
    .B2(net473),
    .X(_0251_));
 sky130_fd_sc_hd__a22o_1 _0940_ (.A1(net477),
    .A2(net407),
    .B1(net398),
    .B2(net484),
    .X(_0252_));
 sky130_fd_sc_hd__or2_1 _0941_ (.A(net87),
    .B(net84),
    .X(_0253_));
 sky130_fd_sc_hd__or4_1 _0942_ (.A(net88),
    .B(net87),
    .C(net85),
    .D(net83),
    .X(_0254_));
 sky130_fd_sc_hd__a22o_1 _0943_ (.A1(net485),
    .A2(net393),
    .B1(net387),
    .B2(net478),
    .X(_0255_));
 sky130_fd_sc_hd__a22o_1 _0944_ (.A1(net454),
    .A2(net393),
    .B1(net387),
    .B2(net447),
    .X(_0256_));
 sky130_fd_sc_hd__a22o_1 _0945_ (.A1(net473),
    .A2(net397),
    .B1(net391),
    .B2(net465),
    .X(_0257_));
 sky130_fd_sc_hd__or2_1 _0946_ (.A(net81),
    .B(net77),
    .X(_0258_));
 sky130_fd_sc_hd__or2_1 _0947_ (.A(net79),
    .B(net59),
    .X(_0259_));
 sky130_fd_sc_hd__a22o_1 _0948_ (.A1(net429),
    .A2(net425),
    .B1(net418),
    .B2(net436),
    .X(_0260_));
 sky130_fd_sc_hd__a22o_1 _0949_ (.A1(net447),
    .A2(net427),
    .B1(net419),
    .B2(net454),
    .X(_0261_));
 sky130_fd_sc_hd__a22o_1 _0950_ (.A1(net478),
    .A2(net427),
    .B1(net419),
    .B2(net485),
    .X(_0262_));
 sky130_fd_sc_hd__a22o_1 _0951_ (.A1(net463),
    .A2(net426),
    .B1(net419),
    .B2(net470),
    .X(_0263_));
 sky130_fd_sc_hd__or2_1 _0952_ (.A(net67),
    .B(net64),
    .X(_0264_));
 sky130_fd_sc_hd__or2_1 _0953_ (.A(net75),
    .B(net68),
    .X(_0265_));
 sky130_fd_sc_hd__or4_2 _0954_ (.A(net75),
    .B(net70),
    .C(net67),
    .D(net65),
    .X(_0266_));
 sky130_fd_sc_hd__or4_1 _0955_ (.A(net217),
    .B(net214),
    .C(_0136_),
    .D(net79),
    .X(_0267_));
 sky130_fd_sc_hd__or4_1 _0956_ (.A(_0133_),
    .B(net211),
    .C(net81),
    .D(net77),
    .X(_0268_));
 sky130_fd_sc_hd__or2_1 _0957_ (.A(net282),
    .B(net208),
    .X(_0269_));
 sky130_fd_sc_hd__or4_1 _0958_ (.A(net287),
    .B(net285),
    .C(net282),
    .D(net208),
    .X(_0270_));
 sky130_fd_sc_hd__or4_1 _0959_ (.A(_0081_),
    .B(_0115_),
    .C(_0130_),
    .D(_0247_),
    .X(_0271_));
 sky130_fd_sc_hd__or4_1 _0960_ (.A(_0090_),
    .B(_0097_),
    .C(_0267_),
    .D(_0268_),
    .X(_0272_));
 sky130_fd_sc_hd__or4_1 _0961_ (.A(_0142_),
    .B(_0225_),
    .C(_0232_),
    .D(_0254_),
    .X(_0273_));
 sky130_fd_sc_hd__or4_1 _0962_ (.A(_0061_),
    .B(_0149_),
    .C(_0266_),
    .D(_0270_),
    .X(_0274_));
 sky130_fd_sc_hd__or4_1 _0963_ (.A(_0051_),
    .B(_0272_),
    .C(_0273_),
    .D(_0274_),
    .X(_0275_));
 sky130_fd_sc_hd__o31a_1 _0964_ (.A1(_0218_),
    .A2(_0271_),
    .A3(_0275_),
    .B1(cs0_reg),
    .X(_0276_));
 sky130_fd_sc_hd__or3_2 _0965_ (.A(net130),
    .B(net128),
    .C(net126),
    .X(_0277_));
 sky130_fd_sc_hd__or2_1 _0966_ (.A(_0164_),
    .B(_0277_),
    .X(_0278_));
 sky130_fd_sc_hd__or2_1 _0967_ (.A(net285),
    .B(net208),
    .X(_0279_));
 sky130_fd_sc_hd__or2_1 _0968_ (.A(net195),
    .B(net193),
    .X(_0280_));
 sky130_fd_sc_hd__or2_1 _0969_ (.A(net278),
    .B(net272),
    .X(_0281_));
 sky130_fd_sc_hd__or2_1 _0970_ (.A(net216),
    .B(net203),
    .X(_0282_));
 sky130_fd_sc_hd__or3_1 _0971_ (.A(_0198_),
    .B(_0204_),
    .C(net135),
    .X(_0283_));
 sky130_fd_sc_hd__or4_1 _0972_ (.A(net145),
    .B(_0198_),
    .C(_0204_),
    .D(net134),
    .X(_0284_));
 sky130_fd_sc_hd__or2_1 _0973_ (.A(net61),
    .B(net207),
    .X(_0285_));
 sky130_fd_sc_hd__or2_1 _0974_ (.A(_0041_),
    .B(net59),
    .X(_0286_));
 sky130_fd_sc_hd__or4_1 _0975_ (.A(net315),
    .B(net313),
    .C(net107),
    .D(net106),
    .X(_0287_));
 sky130_fd_sc_hd__or3_1 _0976_ (.A(net243),
    .B(net240),
    .C(net238),
    .X(_0288_));
 sky130_fd_sc_hd__or4_1 _0977_ (.A(_0285_),
    .B(_0286_),
    .C(_0287_),
    .D(_0288_),
    .X(_0289_));
 sky130_fd_sc_hd__or4_1 _0978_ (.A(net333),
    .B(net288),
    .C(net148),
    .D(net125),
    .X(_0290_));
 sky130_fd_sc_hd__or4_1 _0979_ (.A(net311),
    .B(net98),
    .C(net94),
    .D(_0290_),
    .X(_0291_));
 sky130_fd_sc_hd__or4_1 _0980_ (.A(net294),
    .B(net248),
    .C(net231),
    .D(net225),
    .X(_0292_));
 sky130_fd_sc_hd__or4_1 _0981_ (.A(_0088_),
    .B(_0093_),
    .C(_0291_),
    .D(_0292_),
    .X(_0293_));
 sky130_fd_sc_hd__or4_1 _0982_ (.A(_0180_),
    .B(_0279_),
    .C(_0280_),
    .D(_0281_),
    .X(_0294_));
 sky130_fd_sc_hd__or4_1 _0983_ (.A(net187),
    .B(net183),
    .C(net173),
    .D(net168),
    .X(_0295_));
 sky130_fd_sc_hd__or4_1 _0984_ (.A(net246),
    .B(net120),
    .C(_0282_),
    .D(_0295_),
    .X(_0296_));
 sky130_fd_sc_hd__or4_1 _0985_ (.A(_0278_),
    .B(_0284_),
    .C(_0294_),
    .D(_0296_),
    .X(_0297_));
 sky130_fd_sc_hd__or3_1 _0986_ (.A(_0289_),
    .B(_0293_),
    .C(_0297_),
    .X(_0298_));
 sky130_fd_sc_hd__a22o_1 _0987_ (.A1(net629),
    .A2(net547),
    .B1(net47),
    .B2(_0298_),
    .X(_0000_));
 sky130_fd_sc_hd__or4_2 _0988_ (.A(net313),
    .B(_0031_),
    .C(_0221_),
    .D(net119),
    .X(_0299_));
 sky130_fd_sc_hd__or3_1 _0989_ (.A(net160),
    .B(net157),
    .C(net154),
    .X(_0300_));
 sky130_fd_sc_hd__or2_1 _0990_ (.A(_0677_),
    .B(_0300_),
    .X(_0301_));
 sky130_fd_sc_hd__or3_1 _0991_ (.A(_0056_),
    .B(net206),
    .C(net205),
    .X(_0302_));
 sky130_fd_sc_hd__or3_1 _0992_ (.A(_0059_),
    .B(_0073_),
    .C(_0302_),
    .X(_0303_));
 sky130_fd_sc_hd__or2_1 _0993_ (.A(net240),
    .B(net239),
    .X(_0304_));
 sky130_fd_sc_hd__or3_1 _0994_ (.A(net240),
    .B(net238),
    .C(_0112_),
    .X(_0305_));
 sky130_fd_sc_hd__or4_1 _0995_ (.A(_0243_),
    .B(_0246_),
    .C(_0303_),
    .D(_0305_),
    .X(_0306_));
 sky130_fd_sc_hd__or4_1 _0996_ (.A(net282),
    .B(net268),
    .C(net180),
    .D(net132),
    .X(_0307_));
 sky130_fd_sc_hd__or4_1 _0997_ (.A(net195),
    .B(net191),
    .C(net72),
    .D(net67),
    .X(_0308_));
 sky130_fd_sc_hd__or2_1 _0998_ (.A(_0041_),
    .B(_0169_),
    .X(_0309_));
 sky130_fd_sc_hd__or4_1 _0999_ (.A(_0048_),
    .B(_0089_),
    .C(_0307_),
    .D(_0308_),
    .X(_0310_));
 sky130_fd_sc_hd__or4_1 _1000_ (.A(net253),
    .B(net250),
    .C(net214),
    .D(net103),
    .X(_0311_));
 sky130_fd_sc_hd__or4_1 _1001_ (.A(net228),
    .B(net226),
    .C(net190),
    .D(_0311_),
    .X(_0312_));
 sky130_fd_sc_hd__or4_1 _1002_ (.A(_0277_),
    .B(_0309_),
    .C(_0310_),
    .D(_0312_),
    .X(_0313_));
 sky130_fd_sc_hd__or4_1 _1003_ (.A(_0192_),
    .B(_0199_),
    .C(_0250_),
    .D(net60),
    .X(_0314_));
 sky130_fd_sc_hd__or3_1 _1004_ (.A(_0299_),
    .B(_0301_),
    .C(_0314_),
    .X(_0315_));
 sky130_fd_sc_hd__or3_1 _1005_ (.A(_0306_),
    .B(_0313_),
    .C(_0315_),
    .X(_0316_));
 sky130_fd_sc_hd__a22o_1 _1006_ (.A1(net550),
    .A2(net630),
    .B1(net50),
    .B2(_0316_),
    .X(_0001_));
 sky130_fd_sc_hd__or4_1 _1007_ (.A(net288),
    .B(net225),
    .C(net103),
    .D(net98),
    .X(_0317_));
 sky130_fd_sc_hd__or4_1 _1008_ (.A(_0685_),
    .B(net108),
    .C(net106),
    .D(_0317_),
    .X(_0318_));
 sky130_fd_sc_hd__or4_1 _1009_ (.A(net274),
    .B(net196),
    .C(net175),
    .D(net166),
    .X(_0319_));
 sky130_fd_sc_hd__or4_1 _1010_ (.A(net242),
    .B(net239),
    .C(net218),
    .D(net121),
    .X(_0320_));
 sky130_fd_sc_hd__or4_1 _1011_ (.A(_0050_),
    .B(_0318_),
    .C(_0319_),
    .D(_0320_),
    .X(_0321_));
 sky130_fd_sc_hd__or3_1 _1012_ (.A(_0133_),
    .B(net206),
    .C(net205),
    .X(_0322_));
 sky130_fd_sc_hd__or4_1 _1013_ (.A(net159),
    .B(net157),
    .C(_0209_),
    .D(net126),
    .X(_0323_));
 sky130_fd_sc_hd__or4_1 _1014_ (.A(net212),
    .B(net202),
    .C(net201),
    .D(net82),
    .X(_0324_));
 sky130_fd_sc_hd__or3_1 _1015_ (.A(_0322_),
    .B(_0323_),
    .C(_0324_),
    .X(_0325_));
 sky130_fd_sc_hd__or2_1 _1016_ (.A(net259),
    .B(net252),
    .X(_0326_));
 sky130_fd_sc_hd__or3_1 _1017_ (.A(net258),
    .B(net256),
    .C(net252),
    .X(_0327_));
 sky130_fd_sc_hd__or3_2 _1018_ (.A(net74),
    .B(net71),
    .C(net66),
    .X(_0328_));
 sky130_fd_sc_hd__or2_1 _1019_ (.A(_0327_),
    .B(_0328_),
    .X(_0329_));
 sky130_fd_sc_hd__or2_1 _1020_ (.A(_0190_),
    .B(_0243_),
    .X(_0330_));
 sky130_fd_sc_hd__or3_2 _1021_ (.A(_0073_),
    .B(net89),
    .C(net85),
    .X(_0331_));
 sky130_fd_sc_hd__or4_1 _1022_ (.A(net312),
    .B(net284),
    .C(net267),
    .D(net147),
    .X(_0332_));
 sky130_fd_sc_hd__or3_2 _1023_ (.A(net145),
    .B(net139),
    .C(net136),
    .X(_0333_));
 sky130_fd_sc_hd__or4_1 _1024_ (.A(_0677_),
    .B(net62),
    .C(_0332_),
    .D(_0333_),
    .X(_0334_));
 sky130_fd_sc_hd__or4_1 _1025_ (.A(_0329_),
    .B(_0330_),
    .C(_0331_),
    .D(_0334_),
    .X(_0335_));
 sky130_fd_sc_hd__or3_1 _1026_ (.A(_0321_),
    .B(_0325_),
    .C(_0335_),
    .X(_0336_));
 sky130_fd_sc_hd__a22o_1 _1027_ (.A1(net542),
    .A2(net628),
    .B1(net42),
    .B2(_0336_),
    .X(_0002_));
 sky130_fd_sc_hd__or4_1 _1028_ (.A(net287),
    .B(_0243_),
    .C(net91),
    .D(_0269_),
    .X(_0337_));
 sky130_fd_sc_hd__or4_1 _1029_ (.A(net302),
    .B(net251),
    .C(net244),
    .D(net112),
    .X(_0338_));
 sky130_fd_sc_hd__or2_1 _1030_ (.A(net272),
    .B(net270),
    .X(_0339_));
 sky130_fd_sc_hd__or3_1 _1031_ (.A(net273),
    .B(_0077_),
    .C(net270),
    .X(_0340_));
 sky130_fd_sc_hd__or3_1 _1032_ (.A(net254),
    .B(_0326_),
    .C(_0340_),
    .X(_0341_));
 sky130_fd_sc_hd__or3_1 _1033_ (.A(_0337_),
    .B(_0338_),
    .C(_0341_),
    .X(_0342_));
 sky130_fd_sc_hd__or4_1 _1034_ (.A(net294),
    .B(net292),
    .C(net246),
    .D(net120),
    .X(_0343_));
 sky130_fd_sc_hd__or4_2 _1035_ (.A(_0088_),
    .B(net243),
    .C(net101),
    .D(_0343_),
    .X(_0344_));
 sky130_fd_sc_hd__or4_1 _1036_ (.A(net211),
    .B(net161),
    .C(net142),
    .D(net100),
    .X(_0345_));
 sky130_fd_sc_hd__or2_1 _1037_ (.A(_0171_),
    .B(_0345_),
    .X(_0346_));
 sky130_fd_sc_hd__or2_1 _1038_ (.A(net192),
    .B(net81),
    .X(_0347_));
 sky130_fd_sc_hd__or2_1 _1039_ (.A(net113),
    .B(net104),
    .X(_0348_));
 sky130_fd_sc_hd__or4_1 _1040_ (.A(net70),
    .B(net64),
    .C(_0347_),
    .D(_0348_),
    .X(_0349_));
 sky130_fd_sc_hd__or4_1 _1041_ (.A(net58),
    .B(_0344_),
    .C(_0346_),
    .D(_0349_),
    .X(_0350_));
 sky130_fd_sc_hd__or3_1 _1042_ (.A(net334),
    .B(net332),
    .C(net328),
    .X(_0351_));
 sky130_fd_sc_hd__or4_1 _1043_ (.A(net237),
    .B(net233),
    .C(net181),
    .D(net176),
    .X(_0352_));
 sky130_fd_sc_hd__or3_2 _1044_ (.A(net130),
    .B(net126),
    .C(net124),
    .X(_0353_));
 sky130_fd_sc_hd__or4_1 _1045_ (.A(net223),
    .B(net220),
    .C(net212),
    .D(net204),
    .X(_0354_));
 sky130_fd_sc_hd__or4_1 _1046_ (.A(_0040_),
    .B(_0333_),
    .C(_0353_),
    .D(_0354_),
    .X(_0355_));
 sky130_fd_sc_hd__or4_1 _1047_ (.A(_0074_),
    .B(_0351_),
    .C(_0352_),
    .D(_0355_),
    .X(_0356_));
 sky130_fd_sc_hd__or3_1 _1048_ (.A(_0342_),
    .B(_0350_),
    .C(_0356_),
    .X(_0357_));
 sky130_fd_sc_hd__a22o_1 _1049_ (.A1(net542),
    .A2(net624),
    .B1(net42),
    .B2(_0357_),
    .X(_0003_));
 sky130_fd_sc_hd__or2_1 _1050_ (.A(net305),
    .B(net215),
    .X(_0358_));
 sky130_fd_sc_hd__or4_2 _1051_ (.A(net185),
    .B(net183),
    .C(net114),
    .D(net112),
    .X(_0359_));
 sky130_fd_sc_hd__or2_1 _1052_ (.A(net61),
    .B(_0175_),
    .X(_0360_));
 sky130_fd_sc_hd__or4_1 _1053_ (.A(net242),
    .B(_0114_),
    .C(_0359_),
    .D(_0360_),
    .X(_0361_));
 sky130_fd_sc_hd__or3_1 _1054_ (.A(net333),
    .B(net328),
    .C(net324),
    .X(_0362_));
 sky130_fd_sc_hd__or2_1 _1055_ (.A(net122),
    .B(net118),
    .X(_0363_));
 sky130_fd_sc_hd__or3_1 _1056_ (.A(net121),
    .B(net119),
    .C(net116),
    .X(_0364_));
 sky130_fd_sc_hd__or4_1 _1057_ (.A(net267),
    .B(net263),
    .C(net88),
    .D(net83),
    .X(_0365_));
 sky130_fd_sc_hd__or4_1 _1058_ (.A(_0032_),
    .B(_0362_),
    .C(_0364_),
    .D(_0365_),
    .X(_0366_));
 sky130_fd_sc_hd__or4_1 _1059_ (.A(_0164_),
    .B(_0266_),
    .C(_0341_),
    .D(_0366_),
    .X(_0367_));
 sky130_fd_sc_hd__or4_1 _1060_ (.A(_0064_),
    .B(_0207_),
    .C(_0239_),
    .D(net59),
    .X(_0368_));
 sky130_fd_sc_hd__or3_1 _1061_ (.A(_0041_),
    .B(_0189_),
    .C(_0358_),
    .X(_0369_));
 sky130_fd_sc_hd__or4_1 _1062_ (.A(net290),
    .B(net246),
    .C(net193),
    .D(net125),
    .X(_0370_));
 sky130_fd_sc_hd__or4_1 _1063_ (.A(net170),
    .B(net137),
    .C(net101),
    .D(net94),
    .X(_0371_));
 sky130_fd_sc_hd__or4_1 _1064_ (.A(_0075_),
    .B(net62),
    .C(_0370_),
    .D(_0371_),
    .X(_0372_));
 sky130_fd_sc_hd__or3_1 _1065_ (.A(_0368_),
    .B(_0369_),
    .C(_0372_),
    .X(_0373_));
 sky130_fd_sc_hd__or3_1 _1066_ (.A(_0361_),
    .B(_0367_),
    .C(_0373_),
    .X(_0374_));
 sky130_fd_sc_hd__a22o_1 _1067_ (.A1(net542),
    .A2(net645),
    .B1(net42),
    .B2(_0374_),
    .X(_0004_));
 sky130_fd_sc_hd__or4_2 _1068_ (.A(_0064_),
    .B(net283),
    .C(net61),
    .D(_0139_),
    .X(_0375_));
 sky130_fd_sc_hd__or2_1 _1069_ (.A(_0060_),
    .B(_0238_),
    .X(_0376_));
 sky130_fd_sc_hd__or4_1 _1070_ (.A(net306),
    .B(net297),
    .C(net177),
    .D(net175),
    .X(_0377_));
 sky130_fd_sc_hd__or4_1 _1071_ (.A(net319),
    .B(net315),
    .C(net230),
    .D(_0377_),
    .X(_0378_));
 sky130_fd_sc_hd__or4_1 _1072_ (.A(net277),
    .B(net268),
    .C(net157),
    .D(net154),
    .X(_0379_));
 sky130_fd_sc_hd__or3_1 _1073_ (.A(net94),
    .B(net92),
    .C(_0244_),
    .X(_0380_));
 sky130_fd_sc_hd__or3_1 _1074_ (.A(net217),
    .B(net204),
    .C(net200),
    .X(_0381_));
 sky130_fd_sc_hd__or3_1 _1075_ (.A(net267),
    .B(net262),
    .C(net255),
    .X(_0382_));
 sky130_fd_sc_hd__or4_1 _1076_ (.A(_0107_),
    .B(_0128_),
    .C(_0379_),
    .D(_0382_),
    .X(_0383_));
 sky130_fd_sc_hd__or4_1 _1077_ (.A(_0191_),
    .B(_0328_),
    .C(_0380_),
    .D(_0381_),
    .X(_0384_));
 sky130_fd_sc_hd__or4_1 _1078_ (.A(net167),
    .B(net139),
    .C(net133),
    .D(net128),
    .X(_0385_));
 sky130_fd_sc_hd__or4_1 _1079_ (.A(net236),
    .B(net120),
    .C(net81),
    .D(net80),
    .X(_0386_));
 sky130_fd_sc_hd__or4_1 _1080_ (.A(net331),
    .B(net197),
    .C(net196),
    .D(_0305_),
    .X(_0387_));
 sky130_fd_sc_hd__or4_2 _1081_ (.A(_0384_),
    .B(_0385_),
    .C(_0386_),
    .D(_0387_),
    .X(_0388_));
 sky130_fd_sc_hd__or4_1 _1082_ (.A(net325),
    .B(_0155_),
    .C(_0231_),
    .D(net89),
    .X(_0389_));
 sky130_fd_sc_hd__or4_1 _1083_ (.A(_0375_),
    .B(_0376_),
    .C(_0378_),
    .D(_0389_),
    .X(_0390_));
 sky130_fd_sc_hd__or3_1 _1084_ (.A(_0383_),
    .B(_0388_),
    .C(_0390_),
    .X(_0391_));
 sky130_fd_sc_hd__a22o_1 _1085_ (.A1(net544),
    .A2(net619),
    .B1(net44),
    .B2(_0391_),
    .X(_0005_));
 sky130_fd_sc_hd__or2_1 _1086_ (.A(net248),
    .B(net244),
    .X(_0392_));
 sky130_fd_sc_hd__or2_1 _1087_ (.A(net178),
    .B(net175),
    .X(_0393_));
 sky130_fd_sc_hd__or4_1 _1088_ (.A(net227),
    .B(net220),
    .C(_0392_),
    .D(_0393_),
    .X(_0394_));
 sky130_fd_sc_hd__or4_1 _1089_ (.A(net275),
    .B(net150),
    .C(net90),
    .D(net77),
    .X(_0395_));
 sky130_fd_sc_hd__or4_2 _1090_ (.A(net333),
    .B(net197),
    .C(net72),
    .D(_0395_),
    .X(_0396_));
 sky130_fd_sc_hd__or4_1 _1091_ (.A(net293),
    .B(net291),
    .C(net231),
    .D(net228),
    .X(_0397_));
 sky130_fd_sc_hd__or3_1 _1092_ (.A(net189),
    .B(net184),
    .C(net182),
    .X(_0398_));
 sky130_fd_sc_hd__or4_1 _1093_ (.A(net322),
    .B(net134),
    .C(net112),
    .D(_0398_),
    .X(_0399_));
 sky130_fd_sc_hd__or4_1 _1094_ (.A(net311),
    .B(net307),
    .C(net138),
    .D(net107),
    .X(_0400_));
 sky130_fd_sc_hd__or4_1 _1095_ (.A(_0221_),
    .B(_0237_),
    .C(_0399_),
    .D(_0400_),
    .X(_0401_));
 sky130_fd_sc_hd__or4_1 _1096_ (.A(net172),
    .B(net167),
    .C(net159),
    .D(net155),
    .X(_0402_));
 sky130_fd_sc_hd__or3_1 _1097_ (.A(net88),
    .B(net86),
    .C(net83),
    .X(_0403_));
 sky130_fd_sc_hd__or4_1 _1098_ (.A(net300),
    .B(net296),
    .C(net215),
    .D(net212),
    .X(_0404_));
 sky130_fd_sc_hd__or3_1 _1099_ (.A(_0397_),
    .B(_0402_),
    .C(_0403_),
    .X(_0405_));
 sky130_fd_sc_hd__or4_1 _1100_ (.A(_0200_),
    .B(_0307_),
    .C(_0353_),
    .D(_0404_),
    .X(_0406_));
 sky130_fd_sc_hd__or3_1 _1101_ (.A(_0394_),
    .B(_0396_),
    .C(_0406_),
    .X(_0407_));
 sky130_fd_sc_hd__or3_1 _1102_ (.A(_0401_),
    .B(_0405_),
    .C(_0407_),
    .X(_0408_));
 sky130_fd_sc_hd__a22o_1 _1103_ (.A1(net542),
    .A2(net616),
    .B1(net42),
    .B2(_0408_),
    .X(_0006_));
 sky130_fd_sc_hd__or4_1 _1104_ (.A(net101),
    .B(net95),
    .C(net93),
    .D(net91),
    .X(_0409_));
 sky130_fd_sc_hd__or2_1 _1105_ (.A(net295),
    .B(net287),
    .X(_0410_));
 sky130_fd_sc_hd__or3_1 _1106_ (.A(net215),
    .B(net213),
    .C(net202),
    .X(_0411_));
 sky130_fd_sc_hd__or4_1 _1107_ (.A(net241),
    .B(net239),
    .C(net87),
    .D(net85),
    .X(_0412_));
 sky130_fd_sc_hd__or4_1 _1108_ (.A(net205),
    .B(net186),
    .C(net105),
    .D(net78),
    .X(_0413_));
 sky130_fd_sc_hd__or2_1 _1109_ (.A(_0042_),
    .B(net62),
    .X(_0414_));
 sky130_fd_sc_hd__or4_1 _1110_ (.A(net278),
    .B(net276),
    .C(net180),
    .D(net176),
    .X(_0415_));
 sky130_fd_sc_hd__or3_2 _1111_ (.A(net171),
    .B(net168),
    .C(net164),
    .X(_0416_));
 sky130_fd_sc_hd__or4_1 _1112_ (.A(net318),
    .B(net313),
    .C(net305),
    .D(net301),
    .X(_0417_));
 sky130_fd_sc_hd__or4_1 _1113_ (.A(_0308_),
    .B(_0382_),
    .C(_0416_),
    .D(_0417_),
    .X(_0418_));
 sky130_fd_sc_hd__or4_1 _1114_ (.A(net220),
    .B(net218),
    .C(_0192_),
    .D(_0224_),
    .X(_0419_));
 sky130_fd_sc_hd__or4_1 _1115_ (.A(_0208_),
    .B(_0214_),
    .C(_0413_),
    .D(_0419_),
    .X(_0420_));
 sky130_fd_sc_hd__or4_1 _1116_ (.A(_0409_),
    .B(_0411_),
    .C(_0412_),
    .D(_0415_),
    .X(_0421_));
 sky130_fd_sc_hd__or3_1 _1117_ (.A(_0198_),
    .B(_0392_),
    .C(_0410_),
    .X(_0422_));
 sky130_fd_sc_hd__or4_1 _1118_ (.A(_0301_),
    .B(_0414_),
    .C(_0421_),
    .D(_0422_),
    .X(_0423_));
 sky130_fd_sc_hd__or3_1 _1119_ (.A(_0418_),
    .B(_0420_),
    .C(_0423_),
    .X(_0424_));
 sky130_fd_sc_hd__a22o_1 _1120_ (.A1(net553),
    .A2(net627),
    .B1(net53),
    .B2(_0424_),
    .X(_0007_));
 sky130_fd_sc_hd__or3_1 _1121_ (.A(net250),
    .B(net249),
    .C(net244),
    .X(_0425_));
 sky130_fd_sc_hd__or3_1 _1122_ (.A(net89),
    .B(_0249_),
    .C(_0252_),
    .X(_0426_));
 sky130_fd_sc_hd__or2_1 _1123_ (.A(_0425_),
    .B(_0426_),
    .X(_0427_));
 sky130_fd_sc_hd__or2_1 _1124_ (.A(_0032_),
    .B(_0036_),
    .X(_0428_));
 sky130_fd_sc_hd__or2_1 _1125_ (.A(net139),
    .B(net125),
    .X(_0429_));
 sky130_fd_sc_hd__or4_1 _1126_ (.A(_0133_),
    .B(net199),
    .C(net192),
    .D(net161),
    .X(_0430_));
 sky130_fd_sc_hd__or4_1 _1127_ (.A(net331),
    .B(net271),
    .C(net98),
    .D(net96),
    .X(_0431_));
 sky130_fd_sc_hd__or4_1 _1128_ (.A(net173),
    .B(net168),
    .C(net162),
    .D(net156),
    .X(_0432_));
 sky130_fd_sc_hd__or4_1 _1129_ (.A(_0397_),
    .B(_0415_),
    .C(_0431_),
    .D(_0432_),
    .X(_0433_));
 sky130_fd_sc_hd__or4_1 _1130_ (.A(net270),
    .B(net233),
    .C(net226),
    .D(net144),
    .X(_0434_));
 sky130_fd_sc_hd__or4_1 _1131_ (.A(_0328_),
    .B(_0398_),
    .C(_0430_),
    .D(_0434_),
    .X(_0435_));
 sky130_fd_sc_hd__or4_1 _1132_ (.A(net306),
    .B(net299),
    .C(net92),
    .D(net90),
    .X(_0436_));
 sky130_fd_sc_hd__or3_1 _1133_ (.A(_0114_),
    .B(_0429_),
    .C(_0436_),
    .X(_0437_));
 sky130_fd_sc_hd__or4_1 _1134_ (.A(net333),
    .B(net326),
    .C(net266),
    .D(net264),
    .X(_0438_));
 sky130_fd_sc_hd__or3_1 _1135_ (.A(net59),
    .B(_0326_),
    .C(_0438_),
    .X(_0439_));
 sky130_fd_sc_hd__or4_1 _1136_ (.A(_0433_),
    .B(_0435_),
    .C(_0437_),
    .D(_0439_),
    .X(_0440_));
 sky130_fd_sc_hd__or4_1 _1137_ (.A(net58),
    .B(_0208_),
    .C(_0225_),
    .D(_0232_),
    .X(_0441_));
 sky130_fd_sc_hd__or4_1 _1138_ (.A(_0427_),
    .B(_0428_),
    .C(_0440_),
    .D(_0441_),
    .X(_0442_));
 sky130_fd_sc_hd__a22o_1 _1139_ (.A1(net543),
    .A2(net626),
    .B1(net43),
    .B2(_0442_),
    .X(_0008_));
 sky130_fd_sc_hd__or4_2 _1140_ (.A(net151),
    .B(net149),
    .C(net121),
    .D(net116),
    .X(_0443_));
 sky130_fd_sc_hd__or2_1 _1141_ (.A(net286),
    .B(net283),
    .X(_0444_));
 sky130_fd_sc_hd__or4_1 _1142_ (.A(_0040_),
    .B(_0200_),
    .C(_0381_),
    .D(_0416_),
    .X(_0445_));
 sky130_fd_sc_hd__or4_1 _1143_ (.A(net224),
    .B(net222),
    .C(net85),
    .D(net84),
    .X(_0446_));
 sky130_fd_sc_hd__or4_1 _1144_ (.A(net293),
    .B(net289),
    .C(net71),
    .D(net64),
    .X(_0447_));
 sky130_fd_sc_hd__or2_1 _1145_ (.A(net207),
    .B(net186),
    .X(_0448_));
 sky130_fd_sc_hd__or4_1 _1146_ (.A(net206),
    .B(net186),
    .C(net162),
    .D(net156),
    .X(_0449_));
 sky130_fd_sc_hd__or4_1 _1147_ (.A(net315),
    .B(net260),
    .C(net252),
    .D(net236),
    .X(_0450_));
 sky130_fd_sc_hd__or4_1 _1148_ (.A(net275),
    .B(net107),
    .C(net92),
    .D(_0450_),
    .X(_0451_));
 sky130_fd_sc_hd__or4_1 _1149_ (.A(_0240_),
    .B(_0270_),
    .C(_0445_),
    .D(_0451_),
    .X(_0452_));
 sky130_fd_sc_hd__or4_1 _1150_ (.A(_0259_),
    .B(_0443_),
    .C(_0446_),
    .D(_0447_),
    .X(_0453_));
 sky130_fd_sc_hd__or4_1 _1151_ (.A(_0147_),
    .B(net190),
    .C(net182),
    .D(_0449_),
    .X(_0454_));
 sky130_fd_sc_hd__or4_1 _1152_ (.A(net331),
    .B(net330),
    .C(net135),
    .D(net132),
    .X(_0455_));
 sky130_fd_sc_hd__or4_1 _1153_ (.A(net280),
    .B(net279),
    .C(_0122_),
    .D(_0455_),
    .X(_0456_));
 sky130_fd_sc_hd__or4_1 _1154_ (.A(_0115_),
    .B(_0278_),
    .C(_0454_),
    .D(_0456_),
    .X(_0457_));
 sky130_fd_sc_hd__or3_1 _1155_ (.A(_0452_),
    .B(_0453_),
    .C(_0457_),
    .X(_0458_));
 sky130_fd_sc_hd__a22o_1 _1156_ (.A1(net549),
    .A2(net644),
    .B1(net49),
    .B2(_0458_),
    .X(_0009_));
 sky130_fd_sc_hd__or2_1 _1157_ (.A(net312),
    .B(net310),
    .X(_0459_));
 sky130_fd_sc_hd__or2_1 _1158_ (.A(net280),
    .B(net91),
    .X(_0460_));
 sky130_fd_sc_hd__or4_1 _1159_ (.A(_0098_),
    .B(_0231_),
    .C(_0459_),
    .D(_0460_),
    .X(_0461_));
 sky130_fd_sc_hd__or4_1 _1160_ (.A(net334),
    .B(net327),
    .C(net149),
    .D(net101),
    .X(_0462_));
 sky130_fd_sc_hd__or4_2 _1161_ (.A(net143),
    .B(net139),
    .C(net136),
    .D(net133),
    .X(_0463_));
 sky130_fd_sc_hd__or3_1 _1162_ (.A(net251),
    .B(net248),
    .C(net247),
    .X(_0464_));
 sky130_fd_sc_hd__or4_1 _1163_ (.A(net300),
    .B(net296),
    .C(net121),
    .D(net118),
    .X(_0465_));
 sky130_fd_sc_hd__or4_1 _1164_ (.A(_0462_),
    .B(_0463_),
    .C(_0464_),
    .D(_0465_),
    .X(_0466_));
 sky130_fd_sc_hd__or4_1 _1165_ (.A(net320),
    .B(net223),
    .C(net97),
    .D(net73),
    .X(_0467_));
 sky130_fd_sc_hd__or4_1 _1166_ (.A(_0123_),
    .B(_0171_),
    .C(_0412_),
    .D(_0467_),
    .X(_0468_));
 sky130_fd_sc_hd__or4_1 _1167_ (.A(_0179_),
    .B(_0192_),
    .C(_0339_),
    .D(_0347_),
    .X(_0469_));
 sky130_fd_sc_hd__or4_1 _1168_ (.A(_0058_),
    .B(_0161_),
    .C(_0213_),
    .D(_0282_),
    .X(_0470_));
 sky130_fd_sc_hd__or4_1 _1169_ (.A(_0466_),
    .B(_0468_),
    .C(_0469_),
    .D(_0470_),
    .X(_0471_));
 sky130_fd_sc_hd__or3_1 _1170_ (.A(_0375_),
    .B(_0461_),
    .C(_0471_),
    .X(_0472_));
 sky130_fd_sc_hd__a22o_1 _1171_ (.A1(net548),
    .A2(net640),
    .B1(net48),
    .B2(_0472_),
    .X(_0010_));
 sky130_fd_sc_hd__or2_1 _1172_ (.A(net229),
    .B(net219),
    .X(_0473_));
 sky130_fd_sc_hd__or2_1 _1173_ (.A(_0038_),
    .B(net191),
    .X(_0474_));
 sky130_fd_sc_hd__or2_1 _1174_ (.A(net243),
    .B(net116),
    .X(_0475_));
 sky130_fd_sc_hd__or3_1 _1175_ (.A(net75),
    .B(net68),
    .C(net64),
    .X(_0476_));
 sky130_fd_sc_hd__or4_1 _1176_ (.A(_0189_),
    .B(_0237_),
    .C(_0246_),
    .D(_0280_),
    .X(_0477_));
 sky130_fd_sc_hd__or4_1 _1177_ (.A(_0448_),
    .B(_0473_),
    .C(_0474_),
    .D(_0475_),
    .X(_0478_));
 sky130_fd_sc_hd__or4_1 _1178_ (.A(_0066_),
    .B(_0284_),
    .C(_0477_),
    .D(_0478_),
    .X(_0479_));
 sky130_fd_sc_hd__or3_1 _1179_ (.A(_0230_),
    .B(_0259_),
    .C(_0476_),
    .X(_0480_));
 sky130_fd_sc_hd__or3_1 _1180_ (.A(_0678_),
    .B(_0365_),
    .C(_0417_),
    .X(_0481_));
 sky130_fd_sc_hd__or4_1 _1181_ (.A(net210),
    .B(net176),
    .C(net129),
    .D(net124),
    .X(_0482_));
 sky130_fd_sc_hd__or4_1 _1182_ (.A(_0080_),
    .B(net259),
    .C(net199),
    .D(_0482_),
    .X(_0483_));
 sky130_fd_sc_hd__or3_1 _1183_ (.A(_0075_),
    .B(_0103_),
    .C(_0113_),
    .X(_0484_));
 sky130_fd_sc_hd__or4_1 _1184_ (.A(_0309_),
    .B(_0481_),
    .C(_0483_),
    .D(_0484_),
    .X(_0485_));
 sky130_fd_sc_hd__or3_1 _1185_ (.A(_0479_),
    .B(_0480_),
    .C(_0485_),
    .X(_0486_));
 sky130_fd_sc_hd__a22o_1 _1186_ (.A1(net550),
    .A2(net631),
    .B1(net50),
    .B2(_0486_),
    .X(_0011_));
 sky130_fd_sc_hd__or4_1 _1187_ (.A(net180),
    .B(net178),
    .C(_0194_),
    .D(net142),
    .X(_0487_));
 sky130_fd_sc_hd__or3_2 _1188_ (.A(net231),
    .B(net225),
    .C(net223),
    .X(_0488_));
 sky130_fd_sc_hd__or4_1 _1189_ (.A(net326),
    .B(net88),
    .C(net80),
    .D(net77),
    .X(_0489_));
 sky130_fd_sc_hd__or4_1 _1190_ (.A(net264),
    .B(net261),
    .C(net256),
    .D(net253),
    .X(_0490_));
 sky130_fd_sc_hd__or4_1 _1191_ (.A(net213),
    .B(net200),
    .C(net171),
    .D(net164),
    .X(_0491_));
 sky130_fd_sc_hd__or4_1 _1192_ (.A(net291),
    .B(net281),
    .C(_0162_),
    .D(net146),
    .X(_0492_));
 sky130_fd_sc_hd__or4_1 _1193_ (.A(net285),
    .B(_0288_),
    .C(_0353_),
    .D(_0492_),
    .X(_0493_));
 sky130_fd_sc_hd__or4_1 _1194_ (.A(_0103_),
    .B(net234),
    .C(_0488_),
    .D(_0489_),
    .X(_0494_));
 sky130_fd_sc_hd__or4_1 _1195_ (.A(_0047_),
    .B(_0149_),
    .C(_0493_),
    .D(_0494_),
    .X(_0495_));
 sky130_fd_sc_hd__or3_1 _1196_ (.A(_0487_),
    .B(_0490_),
    .C(_0491_),
    .X(_0496_));
 sky130_fd_sc_hd__or4_1 _1197_ (.A(_0340_),
    .B(_0360_),
    .C(_0476_),
    .D(_0496_),
    .X(_0497_));
 sky130_fd_sc_hd__or4_1 _1198_ (.A(_0380_),
    .B(_0401_),
    .C(_0495_),
    .D(_0497_),
    .X(_0498_));
 sky130_fd_sc_hd__a22o_1 _1199_ (.A1(net547),
    .A2(net637),
    .B1(net47),
    .B2(_0498_),
    .X(_0012_));
 sky130_fd_sc_hd__or2_1 _1200_ (.A(_0157_),
    .B(net181),
    .X(_0499_));
 sky130_fd_sc_hd__or4_1 _1201_ (.A(net297),
    .B(net271),
    .C(net123),
    .D(net115),
    .X(_0500_));
 sky130_fd_sc_hd__or2_1 _1202_ (.A(net261),
    .B(net192),
    .X(_0501_));
 sky130_fd_sc_hd__or4_1 _1203_ (.A(net286),
    .B(net210),
    .C(net152),
    .D(net129),
    .X(_0502_));
 sky130_fd_sc_hd__or4_1 _1204_ (.A(_0107_),
    .B(_0402_),
    .C(_0426_),
    .D(_0443_),
    .X(_0503_));
 sky130_fd_sc_hd__or4_1 _1205_ (.A(_0042_),
    .B(_0238_),
    .C(_0354_),
    .D(_0500_),
    .X(_0504_));
 sky130_fd_sc_hd__or4_1 _1206_ (.A(net74),
    .B(net70),
    .C(_0501_),
    .D(_0502_),
    .X(_0505_));
 sky130_fd_sc_hd__or4_1 _1207_ (.A(_0080_),
    .B(_0096_),
    .C(_0122_),
    .D(net60),
    .X(_0506_));
 sky130_fd_sc_hd__or4_1 _1208_ (.A(_0503_),
    .B(_0504_),
    .C(_0505_),
    .D(_0506_),
    .X(_0507_));
 sky130_fd_sc_hd__or4_1 _1209_ (.A(_0283_),
    .B(_0306_),
    .C(_0499_),
    .D(_0507_),
    .X(_0508_));
 sky130_fd_sc_hd__a22o_1 _1210_ (.A1(net550),
    .A2(net622),
    .B1(net50),
    .B2(_0508_),
    .X(_0013_));
 sky130_fd_sc_hd__or2_1 _1211_ (.A(net137),
    .B(net132),
    .X(_0509_));
 sky130_fd_sc_hd__or4_1 _1212_ (.A(_0148_),
    .B(_0304_),
    .C(_0444_),
    .D(_0509_),
    .X(_0510_));
 sky130_fd_sc_hd__or4_1 _1213_ (.A(_0058_),
    .B(_0073_),
    .C(_0170_),
    .D(_0264_),
    .X(_0511_));
 sky130_fd_sc_hd__or4_1 _1214_ (.A(_0378_),
    .B(_0427_),
    .C(_0510_),
    .D(_0511_),
    .X(_0512_));
 sky130_fd_sc_hd__or3_1 _1215_ (.A(net262),
    .B(net257),
    .C(net254),
    .X(_0513_));
 sky130_fd_sc_hd__or3_1 _1216_ (.A(_0364_),
    .B(_0462_),
    .C(_0513_),
    .X(_0514_));
 sky130_fd_sc_hd__or3_1 _1217_ (.A(net265),
    .B(net153),
    .C(net145),
    .X(_0515_));
 sky130_fd_sc_hd__or4_1 _1218_ (.A(net233),
    .B(net113),
    .C(_0246_),
    .D(_0515_),
    .X(_0516_));
 sky130_fd_sc_hd__or4_1 _1219_ (.A(_0040_),
    .B(_0157_),
    .C(_0514_),
    .D(_0516_),
    .X(_0517_));
 sky130_fd_sc_hd__or3_1 _1220_ (.A(_0325_),
    .B(_0512_),
    .C(_0517_),
    .X(_0518_));
 sky130_fd_sc_hd__a22o_1 _1221_ (.A1(net550),
    .A2(net621),
    .B1(net50),
    .B2(_0518_),
    .X(_0014_));
 sky130_fd_sc_hd__or2_1 _1222_ (.A(_0032_),
    .B(_0403_),
    .X(_0519_));
 sky130_fd_sc_hd__or2_1 _1223_ (.A(net296),
    .B(net82),
    .X(_0520_));
 sky130_fd_sc_hd__or2_1 _1224_ (.A(net308),
    .B(_0112_),
    .X(_0521_));
 sky130_fd_sc_hd__or3_1 _1225_ (.A(net94),
    .B(net91),
    .C(net72),
    .X(_0522_));
 sky130_fd_sc_hd__or4_1 _1226_ (.A(net229),
    .B(net173),
    .C(_0197_),
    .D(net128),
    .X(_0523_));
 sky130_fd_sc_hd__or4_1 _1227_ (.A(net289),
    .B(net111),
    .C(net104),
    .D(net100),
    .X(_0524_));
 sky130_fd_sc_hd__or2_1 _1228_ (.A(_0523_),
    .B(_0524_),
    .X(_0525_));
 sky130_fd_sc_hd__or4_1 _1229_ (.A(net61),
    .B(_0190_),
    .C(net138),
    .D(net135),
    .X(_0526_));
 sky130_fd_sc_hd__or3_1 _1230_ (.A(net197),
    .B(net71),
    .C(net69),
    .X(_0527_));
 sky130_fd_sc_hd__or4_1 _1231_ (.A(_0129_),
    .B(_0513_),
    .C(_0522_),
    .D(_0527_),
    .X(_0528_));
 sky130_fd_sc_hd__or4_1 _1232_ (.A(_0281_),
    .B(_0525_),
    .C(_0526_),
    .D(_0528_),
    .X(_0529_));
 sky130_fd_sc_hd__or4_1 _1233_ (.A(net251),
    .B(net244),
    .C(net237),
    .D(net235),
    .X(_0530_));
 sky130_fd_sc_hd__or4_1 _1234_ (.A(net212),
    .B(net204),
    .C(_0181_),
    .D(_0530_),
    .X(_0531_));
 sky130_fd_sc_hd__or4_1 _1235_ (.A(_0475_),
    .B(_0520_),
    .C(_0521_),
    .D(_0531_),
    .X(_0532_));
 sky130_fd_sc_hd__or4_1 _1236_ (.A(_0499_),
    .B(_0519_),
    .C(_0529_),
    .D(_0532_),
    .X(_0533_));
 sky130_fd_sc_hd__a22o_1 _1237_ (.A1(net543),
    .A2(net632),
    .B1(net43),
    .B2(_0533_),
    .X(_0015_));
 sky130_fd_sc_hd__or3_1 _1238_ (.A(net294),
    .B(net292),
    .C(net290),
    .X(_0534_));
 sky130_fd_sc_hd__or4_1 _1239_ (.A(net321),
    .B(net313),
    .C(net92),
    .D(_0534_),
    .X(_0535_));
 sky130_fd_sc_hd__or2_1 _1240_ (.A(net330),
    .B(net177),
    .X(_0536_));
 sky130_fd_sc_hd__or2_1 _1241_ (.A(net148),
    .B(_0244_),
    .X(_0537_));
 sky130_fd_sc_hd__or3_1 _1242_ (.A(net103),
    .B(net99),
    .C(_0392_),
    .X(_0538_));
 sky130_fd_sc_hd__or3_1 _1243_ (.A(net273),
    .B(_0078_),
    .C(net268),
    .X(_0539_));
 sky130_fd_sc_hd__or4_1 _1244_ (.A(net265),
    .B(net261),
    .C(net129),
    .D(_0210_),
    .X(_0540_));
 sky130_fd_sc_hd__or4_1 _1245_ (.A(_0465_),
    .B(_0476_),
    .C(_0488_),
    .D(_0539_),
    .X(_0541_));
 sky130_fd_sc_hd__or4_1 _1246_ (.A(net209),
    .B(net188),
    .C(net158),
    .D(net144),
    .X(_0542_));
 sky130_fd_sc_hd__or3_1 _1247_ (.A(net279),
    .B(net276),
    .C(net90),
    .X(_0543_));
 sky130_fd_sc_hd__or4_1 _1248_ (.A(_0327_),
    .B(_0432_),
    .C(_0542_),
    .D(_0543_),
    .X(_0544_));
 sky130_fd_sc_hd__or4_1 _1249_ (.A(_0535_),
    .B(_0538_),
    .C(_0541_),
    .D(_0544_),
    .X(_0545_));
 sky130_fd_sc_hd__or4_1 _1250_ (.A(net286),
    .B(net210),
    .C(_0253_),
    .D(_0536_),
    .X(_0546_));
 sky130_fd_sc_hd__or4_1 _1251_ (.A(net137),
    .B(net113),
    .C(net110),
    .D(net104),
    .X(_0547_));
 sky130_fd_sc_hd__or4_1 _1252_ (.A(_0147_),
    .B(net79),
    .C(net78),
    .D(_0547_),
    .X(_0548_));
 sky130_fd_sc_hd__or4_1 _1253_ (.A(_0062_),
    .B(net202),
    .C(_0459_),
    .D(_0540_),
    .X(_0549_));
 sky130_fd_sc_hd__or4_1 _1254_ (.A(_0537_),
    .B(_0546_),
    .C(_0548_),
    .D(_0549_),
    .X(_0550_));
 sky130_fd_sc_hd__or2_1 _1255_ (.A(_0545_),
    .B(_0550_),
    .X(_0551_));
 sky130_fd_sc_hd__a22o_1 _1256_ (.A1(net548),
    .A2(net638),
    .B1(net48),
    .B2(_0551_),
    .X(_0016_));
 sky130_fd_sc_hd__or2_1 _1257_ (.A(net209),
    .B(_0149_),
    .X(_0552_));
 sky130_fd_sc_hd__or2_1 _1258_ (.A(net63),
    .B(net86),
    .X(_0553_));
 sky130_fd_sc_hd__or2_1 _1259_ (.A(net257),
    .B(_0096_),
    .X(_0554_));
 sky130_fd_sc_hd__or2_1 _1260_ (.A(net131),
    .B(_0215_),
    .X(_0555_));
 sky130_fd_sc_hd__or4_1 _1261_ (.A(_0464_),
    .B(_0553_),
    .C(_0554_),
    .D(_0555_),
    .X(_0556_));
 sky130_fd_sc_hd__or4_1 _1262_ (.A(_0040_),
    .B(_0201_),
    .C(_0362_),
    .D(_0447_),
    .X(_0557_));
 sky130_fd_sc_hd__or4_1 _1263_ (.A(net269),
    .B(net100),
    .C(_0250_),
    .D(net79),
    .X(_0558_));
 sky130_fd_sc_hd__or4_1 _1264_ (.A(_0031_),
    .B(_0049_),
    .C(_0204_),
    .D(_0282_),
    .X(_0559_));
 sky130_fd_sc_hd__or4_1 _1265_ (.A(_0135_),
    .B(_0557_),
    .C(_0558_),
    .D(_0559_),
    .X(_0560_));
 sky130_fd_sc_hd__or4_1 _1266_ (.A(net185),
    .B(_0181_),
    .C(_0189_),
    .D(net111),
    .X(_0561_));
 sky130_fd_sc_hd__or4_1 _1267_ (.A(_0172_),
    .B(_0473_),
    .C(_0552_),
    .D(_0561_),
    .X(_0562_));
 sky130_fd_sc_hd__or3_1 _1268_ (.A(_0556_),
    .B(_0560_),
    .C(_0562_),
    .X(_0563_));
 sky130_fd_sc_hd__a22o_1 _1269_ (.A1(net553),
    .A2(net646),
    .B1(net53),
    .B2(_0563_),
    .X(_0017_));
 sky130_fd_sc_hd__or3_1 _1270_ (.A(net223),
    .B(net220),
    .C(net218),
    .X(_0564_));
 sky130_fd_sc_hd__or3_1 _1271_ (.A(net242),
    .B(_0114_),
    .C(_0564_),
    .X(_0565_));
 sky130_fd_sc_hd__or2_1 _1272_ (.A(_0322_),
    .B(_0539_),
    .X(_0566_));
 sky130_fd_sc_hd__or2_1 _1273_ (.A(net123),
    .B(net117),
    .X(_0567_));
 sky130_fd_sc_hd__or4_1 _1274_ (.A(net327),
    .B(net324),
    .C(net151),
    .D(net147),
    .X(_0568_));
 sky130_fd_sc_hd__or3_1 _1275_ (.A(_0074_),
    .B(_0464_),
    .C(_0568_),
    .X(_0569_));
 sky130_fd_sc_hd__or4_1 _1276_ (.A(net108),
    .B(net73),
    .C(_0520_),
    .D(_0567_),
    .X(_0570_));
 sky130_fd_sc_hd__or4_1 _1277_ (.A(net259),
    .B(net215),
    .C(net201),
    .D(net83),
    .X(_0571_));
 sky130_fd_sc_hd__or4_1 _1278_ (.A(net262),
    .B(net255),
    .C(_0410_),
    .D(_0571_),
    .X(_0572_));
 sky130_fd_sc_hd__or4_1 _1279_ (.A(net195),
    .B(_0205_),
    .C(net119),
    .D(net95),
    .X(_0573_));
 sky130_fd_sc_hd__or4_1 _1280_ (.A(_0158_),
    .B(_0323_),
    .C(_0333_),
    .D(_0573_),
    .X(_0574_));
 sky130_fd_sc_hd__or4_1 _1281_ (.A(_0569_),
    .B(_0570_),
    .C(_0572_),
    .D(_0574_),
    .X(_0575_));
 sky130_fd_sc_hd__or4_1 _1282_ (.A(_0428_),
    .B(_0565_),
    .C(_0566_),
    .D(_0575_),
    .X(_0576_));
 sky130_fd_sc_hd__a22o_1 _1283_ (.A1(net543),
    .A2(net636),
    .B1(net43),
    .B2(_0576_),
    .X(_0018_));
 sky130_fd_sc_hd__or4_1 _1284_ (.A(_0337_),
    .B(_0376_),
    .C(_0519_),
    .D(_0566_),
    .X(_0577_));
 sky130_fd_sc_hd__or3_1 _1285_ (.A(net330),
    .B(net303),
    .C(net214),
    .X(_0578_));
 sky130_fd_sc_hd__or4_1 _1286_ (.A(net311),
    .B(net307),
    .C(net195),
    .D(net193),
    .X(_0579_));
 sky130_fd_sc_hd__or4_1 _1287_ (.A(_0191_),
    .B(_0488_),
    .C(_0578_),
    .D(_0579_),
    .X(_0580_));
 sky130_fd_sc_hd__or4_1 _1288_ (.A(_0096_),
    .B(_0106_),
    .C(_0161_),
    .D(_0175_),
    .X(_0581_));
 sky130_fd_sc_hd__or4_1 _1289_ (.A(net280),
    .B(net198),
    .C(net126),
    .D(net80),
    .X(_0582_));
 sky130_fd_sc_hd__or4_1 _1290_ (.A(_0110_),
    .B(net234),
    .C(_0219_),
    .D(_0582_),
    .X(_0583_));
 sky130_fd_sc_hd__or2_1 _1291_ (.A(net190),
    .B(net186),
    .X(_0584_));
 sky130_fd_sc_hd__or4_1 _1292_ (.A(_0170_),
    .B(_0231_),
    .C(_0265_),
    .D(_0584_),
    .X(_0585_));
 sky130_fd_sc_hd__or4_1 _1293_ (.A(_0283_),
    .B(_0581_),
    .C(_0583_),
    .D(_0585_),
    .X(_0586_));
 sky130_fd_sc_hd__or3_1 _1294_ (.A(_0577_),
    .B(_0580_),
    .C(_0586_),
    .X(_0587_));
 sky130_fd_sc_hd__a22o_1 _1295_ (.A1(net546),
    .A2(net618),
    .B1(net46),
    .B2(_0587_),
    .X(_0019_));
 sky130_fd_sc_hd__or3_1 _1296_ (.A(net272),
    .B(net271),
    .C(net268),
    .X(_0588_));
 sky130_fd_sc_hd__or3_1 _1297_ (.A(net189),
    .B(net184),
    .C(net158),
    .X(_0589_));
 sky130_fd_sc_hd__or3_1 _1298_ (.A(net238),
    .B(net236),
    .C(net178),
    .X(_0590_));
 sky130_fd_sc_hd__or4_1 _1299_ (.A(_0090_),
    .B(_0201_),
    .C(_0589_),
    .D(_0590_),
    .X(_0591_));
 sky130_fd_sc_hd__or4_1 _1300_ (.A(_0060_),
    .B(_0491_),
    .C(_0588_),
    .D(_0591_),
    .X(_0592_));
 sky130_fd_sc_hd__or4_1 _1301_ (.A(net74),
    .B(net66),
    .C(_0521_),
    .D(_0536_),
    .X(_0593_));
 sky130_fd_sc_hd__or4_1 _1302_ (.A(_0064_),
    .B(_0148_),
    .C(_0326_),
    .D(_0348_),
    .X(_0594_));
 sky130_fd_sc_hd__or4_1 _1303_ (.A(_0299_),
    .B(_0460_),
    .C(_0593_),
    .D(_0594_),
    .X(_0595_));
 sky130_fd_sc_hd__or4_1 _1304_ (.A(net232),
    .B(net226),
    .C(net222),
    .D(net152),
    .X(_0596_));
 sky130_fd_sc_hd__or4_1 _1305_ (.A(net309),
    .B(_0206_),
    .C(_0239_),
    .D(_0596_),
    .X(_0597_));
 sky130_fd_sc_hd__or4_1 _1306_ (.A(_0277_),
    .B(_0285_),
    .C(_0331_),
    .D(_0597_),
    .X(_0598_));
 sky130_fd_sc_hd__or3_1 _1307_ (.A(_0592_),
    .B(_0595_),
    .C(_0598_),
    .X(_0599_));
 sky130_fd_sc_hd__a22o_1 _1308_ (.A1(net548),
    .A2(net639),
    .B1(net48),
    .B2(_0599_),
    .X(_0020_));
 sky130_fd_sc_hd__or2_1 _1309_ (.A(net278),
    .B(_0522_),
    .X(_0600_));
 sky130_fd_sc_hd__or4_1 _1310_ (.A(_0677_),
    .B(_0060_),
    .C(_0157_),
    .D(_0490_),
    .X(_0601_));
 sky130_fd_sc_hd__or4_1 _1311_ (.A(net208),
    .B(net178),
    .C(net170),
    .D(_0244_),
    .X(_0602_));
 sky130_fd_sc_hd__or4_1 _1312_ (.A(net281),
    .B(net279),
    .C(net228),
    .D(net84),
    .X(_0603_));
 sky130_fd_sc_hd__or4_1 _1313_ (.A(_0142_),
    .B(_0287_),
    .C(_0602_),
    .D(_0603_),
    .X(_0604_));
 sky130_fd_sc_hd__or4_1 _1314_ (.A(_0114_),
    .B(net227),
    .C(net224),
    .D(_0339_),
    .X(_0605_));
 sky130_fd_sc_hd__or4_1 _1315_ (.A(_0047_),
    .B(_0148_),
    .C(_0169_),
    .D(_0363_),
    .X(_0606_));
 sky130_fd_sc_hd__or4_1 _1316_ (.A(_0474_),
    .B(_0604_),
    .C(_0605_),
    .D(_0606_),
    .X(_0607_));
 sky130_fd_sc_hd__or4_1 _1317_ (.A(net58),
    .B(_0217_),
    .C(_0277_),
    .D(_0600_),
    .X(_0608_));
 sky130_fd_sc_hd__or3_1 _1318_ (.A(_0601_),
    .B(_0607_),
    .C(_0608_),
    .X(_0609_));
 sky130_fd_sc_hd__a22o_1 _1319_ (.A1(net554),
    .A2(net643),
    .B1(net54),
    .B2(_0609_),
    .X(_0021_));
 sky130_fd_sc_hd__or4_1 _1320_ (.A(_0180_),
    .B(_0199_),
    .C(_0204_),
    .D(_0304_),
    .X(_0610_));
 sky130_fd_sc_hd__or3_1 _1321_ (.A(_0069_),
    .B(net180),
    .C(net67),
    .X(_0611_));
 sky130_fd_sc_hd__or4_1 _1322_ (.A(net217),
    .B(net199),
    .C(net153),
    .D(net129),
    .X(_0612_));
 sky130_fd_sc_hd__or3_1 _1323_ (.A(_0501_),
    .B(_0584_),
    .C(_0612_),
    .X(_0613_));
 sky130_fd_sc_hd__or3_1 _1324_ (.A(net277),
    .B(net168),
    .C(net164),
    .X(_0614_));
 sky130_fd_sc_hd__or4_1 _1325_ (.A(net233),
    .B(net232),
    .C(net150),
    .D(_0614_),
    .X(_0615_));
 sky130_fd_sc_hd__or4_1 _1326_ (.A(_0610_),
    .B(_0611_),
    .C(_0613_),
    .D(_0615_),
    .X(_0616_));
 sky130_fd_sc_hd__or4_1 _1327_ (.A(net326),
    .B(net310),
    .C(net303),
    .D(net266),
    .X(_0617_));
 sky130_fd_sc_hd__or4_1 _1328_ (.A(net322),
    .B(net304),
    .C(_0279_),
    .D(_0617_),
    .X(_0618_));
 sky130_fd_sc_hd__or4_1 _1329_ (.A(_0446_),
    .B(_0535_),
    .C(_0554_),
    .D(_0618_),
    .X(_0619_));
 sky130_fd_sc_hd__or4_1 _1330_ (.A(_0230_),
    .B(_0588_),
    .C(_0616_),
    .D(_0619_),
    .X(_0620_));
 sky130_fd_sc_hd__a22o_1 _1331_ (.A1(net548),
    .A2(net642),
    .B1(net48),
    .B2(_0620_),
    .X(_0022_));
 sky130_fd_sc_hd__or4_1 _1332_ (.A(net189),
    .B(net182),
    .C(net173),
    .D(net164),
    .X(_0621_));
 sky130_fd_sc_hd__or4_2 _1333_ (.A(_0253_),
    .B(net74),
    .C(net66),
    .D(_0621_),
    .X(_0622_));
 sky130_fd_sc_hd__or3_1 _1334_ (.A(_0358_),
    .B(_0393_),
    .C(_0579_),
    .X(_0623_));
 sky130_fd_sc_hd__or2_1 _1335_ (.A(net258),
    .B(net235),
    .X(_0624_));
 sky130_fd_sc_hd__or4_1 _1336_ (.A(_0031_),
    .B(_0224_),
    .C(_0269_),
    .D(_0624_),
    .X(_0625_));
 sky130_fd_sc_hd__or4_1 _1337_ (.A(_0565_),
    .B(_0622_),
    .C(_0623_),
    .D(_0625_),
    .X(_0626_));
 sky130_fd_sc_hd__or4_1 _1338_ (.A(_0379_),
    .B(_0431_),
    .C(_0463_),
    .D(_0555_),
    .X(_0627_));
 sky130_fd_sc_hd__or4_1 _1339_ (.A(net304),
    .B(net294),
    .C(net290),
    .D(net230),
    .X(_0629_));
 sky130_fd_sc_hd__or4_1 _1340_ (.A(_0089_),
    .B(_0330_),
    .C(_0338_),
    .D(_0629_),
    .X(_0630_));
 sky130_fd_sc_hd__or3_1 _1341_ (.A(_0626_),
    .B(_0627_),
    .C(_0630_),
    .X(_0631_));
 sky130_fd_sc_hd__a22o_1 _1342_ (.A1(net547),
    .A2(net634),
    .B1(net47),
    .B2(_0631_),
    .X(_0023_));
 sky130_fd_sc_hd__or4_1 _1343_ (.A(_0041_),
    .B(_0059_),
    .C(net63),
    .D(_0215_),
    .X(_0632_));
 sky130_fd_sc_hd__or3_1 _1344_ (.A(_0685_),
    .B(_0509_),
    .C(_0567_),
    .X(_0633_));
 sky130_fd_sc_hd__or4_1 _1345_ (.A(_0552_),
    .B(_0600_),
    .C(_0632_),
    .D(_0633_),
    .X(_0634_));
 sky130_fd_sc_hd__or3_1 _1346_ (.A(_0488_),
    .B(_0538_),
    .C(_0568_),
    .X(_0635_));
 sky130_fd_sc_hd__or3_1 _1347_ (.A(net262),
    .B(net221),
    .C(net170),
    .X(_0636_));
 sky130_fd_sc_hd__or4_1 _1348_ (.A(_0048_),
    .B(_0300_),
    .C(_0340_),
    .D(_0636_),
    .X(_0637_));
 sky130_fd_sc_hd__or4_1 _1349_ (.A(_0359_),
    .B(_0411_),
    .C(_0426_),
    .D(_0637_),
    .X(_0639_));
 sky130_fd_sc_hd__or4_1 _1350_ (.A(_0487_),
    .B(_0634_),
    .C(_0635_),
    .D(_0639_),
    .X(_0640_));
 sky130_fd_sc_hd__a22o_1 _1351_ (.A1(net544),
    .A2(net617),
    .B1(net44),
    .B2(_0640_),
    .X(_0024_));
 sky130_fd_sc_hd__or3_1 _1352_ (.A(net325),
    .B(net171),
    .C(net169),
    .X(_0641_));
 sky130_fd_sc_hd__or4_1 _1353_ (.A(_0032_),
    .B(_0128_),
    .C(_0352_),
    .D(_0404_),
    .X(_0642_));
 sky130_fd_sc_hd__or4_1 _1354_ (.A(_0409_),
    .B(_0425_),
    .C(_0553_),
    .D(_0641_),
    .X(_0643_));
 sky130_fd_sc_hd__or4_1 _1355_ (.A(net306),
    .B(_0075_),
    .C(net150),
    .D(net134),
    .X(_0644_));
 sky130_fd_sc_hd__or4_1 _1356_ (.A(net310),
    .B(net309),
    .C(net152),
    .D(net146),
    .X(_0645_));
 sky130_fd_sc_hd__or4_1 _1357_ (.A(_0155_),
    .B(net156),
    .C(net122),
    .D(_0645_),
    .X(_0646_));
 sky130_fd_sc_hd__or4_1 _1358_ (.A(_0207_),
    .B(net107),
    .C(net72),
    .D(_0429_),
    .X(_0647_));
 sky130_fd_sc_hd__or4_1 _1359_ (.A(_0066_),
    .B(_0644_),
    .C(_0646_),
    .D(_0647_),
    .X(_0649_));
 sky130_fd_sc_hd__or3_1 _1360_ (.A(_0642_),
    .B(_0643_),
    .C(_0649_),
    .X(_0650_));
 sky130_fd_sc_hd__a22o_1 _1361_ (.A1(net543),
    .A2(net633),
    .B1(net43),
    .B2(_0650_),
    .X(_0025_));
 sky130_fd_sc_hd__or3_1 _1362_ (.A(net216),
    .B(net213),
    .C(_0232_),
    .X(_0651_));
 sky130_fd_sc_hd__or3_1 _1363_ (.A(_0208_),
    .B(_0425_),
    .C(_0651_),
    .X(_0652_));
 sky130_fd_sc_hd__or3_1 _1364_ (.A(net314),
    .B(_0212_),
    .C(net70),
    .X(_0653_));
 sky130_fd_sc_hd__or4_1 _1365_ (.A(net63),
    .B(net177),
    .C(net163),
    .D(_0653_),
    .X(_0654_));
 sky130_fd_sc_hd__or3_1 _1366_ (.A(_0179_),
    .B(_0264_),
    .C(_0537_),
    .X(_0655_));
 sky130_fd_sc_hd__or2_1 _1367_ (.A(_0158_),
    .B(_0240_),
    .X(_0656_));
 sky130_fd_sc_hd__or4_1 _1368_ (.A(_0641_),
    .B(_0654_),
    .C(_0655_),
    .D(_0656_),
    .X(_0657_));
 sky130_fd_sc_hd__or4_1 _1369_ (.A(_0081_),
    .B(_0414_),
    .C(_0652_),
    .D(_0657_),
    .X(_0659_));
 sky130_fd_sc_hd__a22o_1 _1370_ (.A1(net551),
    .A2(net635),
    .B1(net51),
    .B2(_0659_),
    .X(_0026_));
 sky130_fd_sc_hd__or3_1 _1371_ (.A(_0113_),
    .B(_0169_),
    .C(_0254_),
    .X(_0660_));
 sky130_fd_sc_hd__or4_1 _1372_ (.A(_0050_),
    .B(_0158_),
    .C(net58),
    .D(_0351_),
    .X(_0661_));
 sky130_fd_sc_hd__or3_1 _1373_ (.A(_0247_),
    .B(_0278_),
    .C(_0660_),
    .X(_0662_));
 sky130_fd_sc_hd__or3_1 _1374_ (.A(_0652_),
    .B(_0661_),
    .C(_0662_),
    .X(_0663_));
 sky130_fd_sc_hd__a22o_1 _1375_ (.A1(net551),
    .A2(net620),
    .B1(net51),
    .B2(_0663_),
    .X(_0027_));
 sky130_fd_sc_hd__or3_1 _1376_ (.A(net247),
    .B(_0201_),
    .C(_0225_),
    .X(_0664_));
 sky130_fd_sc_hd__or4_1 _1377_ (.A(_0051_),
    .B(_0183_),
    .C(_0651_),
    .D(_0664_),
    .X(_0665_));
 sky130_fd_sc_hd__a22o_1 _1378_ (.A1(net553),
    .A2(net625),
    .B1(net53),
    .B2(_0665_),
    .X(_0028_));
 sky130_fd_sc_hd__or4_1 _1379_ (.A(_0130_),
    .B(net203),
    .C(net201),
    .D(_0218_),
    .X(_0667_));
 sky130_fd_sc_hd__a22o_1 _1380_ (.A1(net553),
    .A2(net623),
    .B1(net53),
    .B2(_0667_),
    .X(_0029_));
 sky130_fd_sc_hd__a21o_1 _1381_ (.A1(net554),
    .A2(net641),
    .B1(net54),
    .X(_0030_));
 sky130_fd_sc_hd__dfxtp_1 _1382_ (.CLK(clknet_2_1__leaf_clk0),
    .D(_0000_),
    .Q(net10));
 sky130_fd_sc_hd__dfxtp_1 _1383_ (.CLK(clknet_2_1__leaf_clk0),
    .D(_0001_),
    .Q(net21));
 sky130_fd_sc_hd__dfxtp_1 _1384_ (.CLK(clknet_2_2__leaf_clk0),
    .D(_0002_),
    .Q(net32));
 sky130_fd_sc_hd__dfxtp_1 _1385_ (.CLK(clknet_2_2__leaf_clk0),
    .D(_0003_),
    .Q(net35));
 sky130_fd_sc_hd__dfxtp_1 _1386_ (.CLK(clknet_2_2__leaf_clk0),
    .D(_0004_),
    .Q(net36));
 sky130_fd_sc_hd__dfxtp_1 _1387_ (.CLK(clknet_2_2__leaf_clk0),
    .D(_0005_),
    .Q(net37));
 sky130_fd_sc_hd__dfxtp_1 _1388_ (.CLK(clknet_2_2__leaf_clk0),
    .D(_0006_),
    .Q(net38));
 sky130_fd_sc_hd__dfxtp_1 _1389_ (.CLK(clknet_2_3__leaf_clk0),
    .D(_0007_),
    .Q(net39));
 sky130_fd_sc_hd__dfxtp_1 _1390_ (.CLK(clknet_2_2__leaf_clk0),
    .D(_0008_),
    .Q(net40));
 sky130_fd_sc_hd__dfxtp_1 _1391_ (.CLK(clknet_2_1__leaf_clk0),
    .D(_0009_),
    .Q(net41));
 sky130_fd_sc_hd__dfxtp_1 _1392_ (.CLK(clknet_2_3__leaf_clk0),
    .D(_0010_),
    .Q(net11));
 sky130_fd_sc_hd__dfxtp_1 _1393_ (.CLK(clknet_2_1__leaf_clk0),
    .D(_0011_),
    .Q(net12));
 sky130_fd_sc_hd__dfxtp_1 _1394_ (.CLK(clknet_2_2__leaf_clk0),
    .D(_0012_),
    .Q(net13));
 sky130_fd_sc_hd__dfxtp_1 _1395_ (.CLK(clknet_2_3__leaf_clk0),
    .D(_0013_),
    .Q(net14));
 sky130_fd_sc_hd__dfxtp_1 _1396_ (.CLK(clknet_2_3__leaf_clk0),
    .D(_0014_),
    .Q(net15));
 sky130_fd_sc_hd__dfxtp_1 _1397_ (.CLK(clknet_2_2__leaf_clk0),
    .D(_0015_),
    .Q(net16));
 sky130_fd_sc_hd__dfxtp_1 _1398_ (.CLK(clknet_2_1__leaf_clk0),
    .D(_0016_),
    .Q(net17));
 sky130_fd_sc_hd__dfxtp_1 _1399_ (.CLK(clknet_2_3__leaf_clk0),
    .D(_0017_),
    .Q(net18));
 sky130_fd_sc_hd__dfxtp_1 _1400_ (.CLK(clknet_2_2__leaf_clk0),
    .D(_0018_),
    .Q(net19));
 sky130_fd_sc_hd__dfxtp_1 _1401_ (.CLK(clknet_2_2__leaf_clk0),
    .D(_0019_),
    .Q(net20));
 sky130_fd_sc_hd__dfxtp_1 _1402_ (.CLK(clknet_2_1__leaf_clk0),
    .D(_0020_),
    .Q(net22));
 sky130_fd_sc_hd__dfxtp_1 _1403_ (.CLK(clknet_2_3__leaf_clk0),
    .D(_0021_),
    .Q(net23));
 sky130_fd_sc_hd__dfxtp_1 _1404_ (.CLK(clknet_2_1__leaf_clk0),
    .D(_0022_),
    .Q(net24));
 sky130_fd_sc_hd__dfxtp_1 _1405_ (.CLK(clknet_2_2__leaf_clk0),
    .D(_0023_),
    .Q(net25));
 sky130_fd_sc_hd__dfxtp_1 _1406_ (.CLK(clknet_2_3__leaf_clk0),
    .D(_0024_),
    .Q(net26));
 sky130_fd_sc_hd__dfxtp_1 _1407_ (.CLK(clknet_2_2__leaf_clk0),
    .D(_0025_),
    .Q(net27));
 sky130_fd_sc_hd__dfxtp_1 _1408_ (.CLK(clknet_2_1__leaf_clk0),
    .D(_0026_),
    .Q(net28));
 sky130_fd_sc_hd__dfxtp_1 _1409_ (.CLK(clknet_2_3__leaf_clk0),
    .D(_0027_),
    .Q(net29));
 sky130_fd_sc_hd__dfxtp_1 _1410_ (.CLK(clknet_2_3__leaf_clk0),
    .D(_0028_),
    .Q(net30));
 sky130_fd_sc_hd__dfxtp_1 _1411_ (.CLK(clknet_2_3__leaf_clk0),
    .D(_0029_),
    .Q(net31));
 sky130_fd_sc_hd__dfxtp_1 _1412_ (.CLK(clknet_2_3__leaf_clk0),
    .D(_0030_),
    .Q(net34));
 sky130_fd_sc_hd__dfxtp_1 _1413_ (.CLK(clknet_2_0__leaf_clk0),
    .D(net1),
    .Q(\addr0_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1414_ (.CLK(clknet_2_0__leaf_clk0),
    .D(net2),
    .Q(\addr0_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1415_ (.CLK(clknet_2_0__leaf_clk0),
    .D(net3),
    .Q(\addr0_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1416_ (.CLK(clknet_2_0__leaf_clk0),
    .D(net4),
    .Q(\addr0_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1417_ (.CLK(clknet_2_0__leaf_clk0),
    .D(net5),
    .Q(\addr0_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1418_ (.CLK(clknet_2_0__leaf_clk0),
    .D(net6),
    .Q(\addr0_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1419_ (.CLK(clknet_2_0__leaf_clk0),
    .D(net7),
    .Q(\addr0_reg[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1420_ (.CLK(clknet_2_0__leaf_clk0),
    .D(net8),
    .Q(\addr0_reg[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1421_ (.CLK(clknet_2_3__leaf_clk0),
    .D(net9),
    .Q(cs0_reg));
 sky130_fd_sc_hd__clkbuf_1 _1422_ (.A(net34),
    .X(net33));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_443 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(addr0[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(addr0[1]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(addr0[2]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(addr0[3]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(addr0[4]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(addr0[5]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(addr0[6]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(addr0[7]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(cs0),
    .X(net9));
 sky130_fd_sc_hd__buf_2 output10 (.A(net10),
    .X(dout0[0]));
 sky130_fd_sc_hd__clkbuf_4 output11 (.A(net11),
    .X(dout0[10]));
 sky130_fd_sc_hd__buf_2 output12 (.A(net12),
    .X(dout0[11]));
 sky130_fd_sc_hd__buf_2 output13 (.A(net13),
    .X(dout0[12]));
 sky130_fd_sc_hd__buf_2 output14 (.A(net14),
    .X(dout0[13]));
 sky130_fd_sc_hd__buf_2 output15 (.A(net15),
    .X(dout0[14]));
 sky130_fd_sc_hd__buf_2 output16 (.A(net16),
    .X(dout0[15]));
 sky130_fd_sc_hd__clkbuf_4 output17 (.A(net17),
    .X(dout0[16]));
 sky130_fd_sc_hd__buf_2 output18 (.A(net18),
    .X(dout0[17]));
 sky130_fd_sc_hd__buf_2 output19 (.A(net19),
    .X(dout0[18]));
 sky130_fd_sc_hd__buf_2 output20 (.A(net20),
    .X(dout0[19]));
 sky130_fd_sc_hd__buf_2 output21 (.A(net21),
    .X(dout0[1]));
 sky130_fd_sc_hd__clkbuf_4 output22 (.A(net22),
    .X(dout0[20]));
 sky130_fd_sc_hd__clkbuf_4 output23 (.A(net23),
    .X(dout0[21]));
 sky130_fd_sc_hd__clkbuf_4 output24 (.A(net24),
    .X(dout0[22]));
 sky130_fd_sc_hd__buf_2 output25 (.A(net25),
    .X(dout0[23]));
 sky130_fd_sc_hd__buf_2 output26 (.A(net26),
    .X(dout0[24]));
 sky130_fd_sc_hd__buf_2 output27 (.A(net27),
    .X(dout0[25]));
 sky130_fd_sc_hd__buf_2 output28 (.A(net28),
    .X(dout0[26]));
 sky130_fd_sc_hd__buf_2 output29 (.A(net29),
    .X(dout0[27]));
 sky130_fd_sc_hd__buf_2 output30 (.A(net30),
    .X(dout0[28]));
 sky130_fd_sc_hd__buf_2 output31 (.A(net31),
    .X(dout0[29]));
 sky130_fd_sc_hd__buf_2 output32 (.A(net32),
    .X(dout0[2]));
 sky130_fd_sc_hd__buf_2 output33 (.A(net33),
    .X(dout0[30]));
 sky130_fd_sc_hd__buf_2 output34 (.A(net34),
    .X(dout0[31]));
 sky130_fd_sc_hd__buf_2 output35 (.A(net35),
    .X(dout0[3]));
 sky130_fd_sc_hd__buf_2 output36 (.A(net36),
    .X(dout0[4]));
 sky130_fd_sc_hd__buf_2 output37 (.A(net37),
    .X(dout0[5]));
 sky130_fd_sc_hd__buf_2 output38 (.A(net38),
    .X(dout0[6]));
 sky130_fd_sc_hd__buf_2 output39 (.A(net39),
    .X(dout0[7]));
 sky130_fd_sc_hd__buf_2 output40 (.A(net40),
    .X(dout0[8]));
 sky130_fd_sc_hd__clkbuf_4 output41 (.A(net41),
    .X(dout0[9]));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout42 (.A(net46),
    .X(net42));
 sky130_fd_sc_hd__buf_1 fanout43 (.A(net45),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 fanout44 (.A(net45),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 fanout45 (.A(net46),
    .X(net45));
 sky130_fd_sc_hd__buf_1 fanout46 (.A(net47),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_2 fanout47 (.A(net57),
    .X(net47));
 sky130_fd_sc_hd__buf_1 fanout48 (.A(net49),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_1 fanout49 (.A(net56),
    .X(net49));
 sky130_fd_sc_hd__buf_1 fanout50 (.A(net52),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 fanout51 (.A(net52),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 fanout52 (.A(net55),
    .X(net52));
 sky130_fd_sc_hd__buf_1 fanout53 (.A(net54),
    .X(net53));
 sky130_fd_sc_hd__buf_1 fanout54 (.A(net55),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 fanout55 (.A(net56),
    .X(net55));
 sky130_fd_sc_hd__buf_1 fanout56 (.A(net57),
    .X(net56));
 sky130_fd_sc_hd__buf_1 fanout57 (.A(_0276_),
    .X(net57));
 sky130_fd_sc_hd__buf_1 fanout58 (.A(_0193_),
    .X(net58));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout59 (.A(_0258_),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 fanout60 (.A(_0258_),
    .X(net60));
 sky130_fd_sc_hd__buf_1 fanout61 (.A(_0135_),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_2 fanout62 (.A(_0123_),
    .X(net62));
 sky130_fd_sc_hd__buf_1 fanout63 (.A(_0110_),
    .X(net63));
 sky130_fd_sc_hd__buf_1 fanout64 (.A(net65),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_1 fanout65 (.A(net66),
    .X(net65));
 sky130_fd_sc_hd__buf_1 fanout66 (.A(_0263_),
    .X(net66));
 sky130_fd_sc_hd__buf_1 fanout67 (.A(net69),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_1 fanout68 (.A(net69),
    .X(net68));
 sky130_fd_sc_hd__buf_1 fanout69 (.A(_0262_),
    .X(net69));
 sky130_fd_sc_hd__buf_1 fanout70 (.A(net71),
    .X(net70));
 sky130_fd_sc_hd__buf_1 fanout71 (.A(_0261_),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_2 fanout72 (.A(net76),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_1 fanout73 (.A(net76),
    .X(net73));
 sky130_fd_sc_hd__buf_1 fanout74 (.A(net76),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_1 fanout75 (.A(net76),
    .X(net75));
 sky130_fd_sc_hd__buf_2 fanout76 (.A(_0260_),
    .X(net76));
 sky130_fd_sc_hd__buf_1 fanout77 (.A(_0257_),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_1 fanout78 (.A(_0257_),
    .X(net78));
 sky130_fd_sc_hd__buf_1 fanout79 (.A(net80),
    .X(net79));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout80 (.A(_0256_),
    .X(net80));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout81 (.A(_0255_),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_1 fanout82 (.A(_0255_),
    .X(net82));
 sky130_fd_sc_hd__buf_1 fanout83 (.A(net84),
    .X(net83));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout84 (.A(_0252_),
    .X(net84));
 sky130_fd_sc_hd__buf_1 fanout85 (.A(_0251_),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_1 fanout86 (.A(_0251_),
    .X(net86));
 sky130_fd_sc_hd__buf_1 fanout87 (.A(_0249_),
    .X(net87));
 sky130_fd_sc_hd__buf_1 fanout88 (.A(_0248_),
    .X(net88));
 sky130_fd_sc_hd__buf_1 fanout89 (.A(_0248_),
    .X(net89));
 sky130_fd_sc_hd__buf_1 fanout90 (.A(_0245_),
    .X(net90));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout91 (.A(_0245_),
    .X(net91));
 sky130_fd_sc_hd__buf_1 fanout92 (.A(_0242_),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_1 fanout93 (.A(_0242_),
    .X(net93));
 sky130_fd_sc_hd__buf_1 fanout94 (.A(_0241_),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_1 fanout95 (.A(_0241_),
    .X(net95));
 sky130_fd_sc_hd__buf_1 fanout96 (.A(_0236_),
    .X(net96));
 sky130_fd_sc_hd__buf_1 fanout97 (.A(_0236_),
    .X(net97));
 sky130_fd_sc_hd__buf_1 fanout98 (.A(net99),
    .X(net98));
 sky130_fd_sc_hd__buf_1 fanout99 (.A(net100),
    .X(net99));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout100 (.A(_0235_),
    .X(net100));
 sky130_fd_sc_hd__buf_1 fanout101 (.A(_0234_),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_1 fanout102 (.A(_0234_),
    .X(net102));
 sky130_fd_sc_hd__buf_1 fanout103 (.A(_0233_),
    .X(net103));
 sky130_fd_sc_hd__buf_1 fanout104 (.A(net106),
    .X(net104));
 sky130_fd_sc_hd__buf_1 fanout105 (.A(net106),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_2 fanout106 (.A(_0229_),
    .X(net106));
 sky130_fd_sc_hd__buf_1 fanout107 (.A(net109),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_1 fanout108 (.A(net109),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_2 fanout109 (.A(_0228_),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_1 fanout110 (.A(_0228_),
    .X(net110));
 sky130_fd_sc_hd__buf_1 fanout111 (.A(net112),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_2 fanout112 (.A(_0227_),
    .X(net112));
 sky130_fd_sc_hd__buf_1 fanout113 (.A(net115),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_1 fanout114 (.A(net115),
    .X(net114));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout115 (.A(_0226_),
    .X(net115));
 sky130_fd_sc_hd__buf_1 fanout116 (.A(net118),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_1 fanout117 (.A(net118),
    .X(net117));
 sky130_fd_sc_hd__buf_1 fanout118 (.A(_0223_),
    .X(net118));
 sky130_fd_sc_hd__buf_1 fanout119 (.A(net120),
    .X(net119));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout120 (.A(_0222_),
    .X(net120));
 sky130_fd_sc_hd__buf_1 fanout121 (.A(net122),
    .X(net121));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout122 (.A(_0220_),
    .X(net122));
 sky130_fd_sc_hd__buf_1 fanout123 (.A(_0219_),
    .X(net123));
 sky130_fd_sc_hd__buf_1 fanout124 (.A(net125),
    .X(net124));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout125 (.A(_0212_),
    .X(net125));
 sky130_fd_sc_hd__buf_1 fanout126 (.A(_0211_),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_1 fanout127 (.A(_0211_),
    .X(net127));
 sky130_fd_sc_hd__buf_1 fanout128 (.A(_0210_),
    .X(net128));
 sky130_fd_sc_hd__buf_1 fanout129 (.A(net131),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_1 fanout130 (.A(net131),
    .X(net130));
 sky130_fd_sc_hd__buf_1 fanout131 (.A(_0209_),
    .X(net131));
 sky130_fd_sc_hd__buf_1 fanout132 (.A(net133),
    .X(net132));
 sky130_fd_sc_hd__buf_1 fanout133 (.A(_0206_),
    .X(net133));
 sky130_fd_sc_hd__buf_1 fanout134 (.A(net135),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_2 fanout135 (.A(_0205_),
    .X(net135));
 sky130_fd_sc_hd__buf_1 fanout136 (.A(_0203_),
    .X(net136));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout137 (.A(net138),
    .X(net137));
 sky130_fd_sc_hd__buf_2 fanout138 (.A(_0202_),
    .X(net138));
 sky130_fd_sc_hd__buf_1 fanout139 (.A(net140),
    .X(net139));
 sky130_fd_sc_hd__buf_1 fanout140 (.A(_0197_),
    .X(net140));
 sky130_fd_sc_hd__buf_1 fanout141 (.A(net142),
    .X(net141));
 sky130_fd_sc_hd__buf_1 fanout142 (.A(net143),
    .X(net142));
 sky130_fd_sc_hd__buf_1 fanout143 (.A(_0196_),
    .X(net143));
 sky130_fd_sc_hd__buf_1 fanout144 (.A(_0195_),
    .X(net144));
 sky130_fd_sc_hd__buf_1 fanout145 (.A(_0194_),
    .X(net145));
 sky130_fd_sc_hd__buf_1 fanout146 (.A(_0188_),
    .X(net146));
 sky130_fd_sc_hd__buf_1 fanout147 (.A(_0188_),
    .X(net147));
 sky130_fd_sc_hd__buf_1 fanout148 (.A(_0187_),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_1 fanout149 (.A(_0187_),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_2 fanout150 (.A(_0186_),
    .X(net150));
 sky130_fd_sc_hd__buf_1 fanout151 (.A(_0186_),
    .X(net151));
 sky130_fd_sc_hd__buf_1 fanout152 (.A(_0185_),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_1 fanout153 (.A(_0185_),
    .X(net153));
 sky130_fd_sc_hd__buf_1 fanout154 (.A(net155),
    .X(net154));
 sky130_fd_sc_hd__buf_1 fanout155 (.A(net156),
    .X(net155));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout156 (.A(_0178_),
    .X(net156));
 sky130_fd_sc_hd__buf_1 fanout157 (.A(net158),
    .X(net157));
 sky130_fd_sc_hd__buf_1 fanout158 (.A(_0176_),
    .X(net158));
 sky130_fd_sc_hd__buf_1 fanout159 (.A(net160),
    .X(net159));
 sky130_fd_sc_hd__buf_1 fanout160 (.A(net161),
    .X(net160));
 sky130_fd_sc_hd__buf_1 fanout161 (.A(_0174_),
    .X(net161));
 sky130_fd_sc_hd__buf_1 fanout162 (.A(_0173_),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_1 fanout163 (.A(_0173_),
    .X(net163));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout164 (.A(net166),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_1 fanout165 (.A(net166),
    .X(net165));
 sky130_fd_sc_hd__buf_1 fanout166 (.A(_0168_),
    .X(net166));
 sky130_fd_sc_hd__clkbuf_2 fanout167 (.A(_0167_),
    .X(net167));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout168 (.A(_0166_),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_1 fanout169 (.A(net170),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_2 fanout170 (.A(_0166_),
    .X(net170));
 sky130_fd_sc_hd__buf_1 fanout171 (.A(net174),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_1 fanout172 (.A(net174),
    .X(net172));
 sky130_fd_sc_hd__buf_1 fanout173 (.A(_0165_),
    .X(net173));
 sky130_fd_sc_hd__buf_1 fanout174 (.A(_0165_),
    .X(net174));
 sky130_fd_sc_hd__buf_1 fanout175 (.A(_0163_),
    .X(net175));
 sky130_fd_sc_hd__buf_1 fanout176 (.A(_0163_),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_2 fanout177 (.A(_0162_),
    .X(net177));
 sky130_fd_sc_hd__buf_1 fanout178 (.A(_0160_),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_1 fanout179 (.A(_0160_),
    .X(net179));
 sky130_fd_sc_hd__buf_1 fanout180 (.A(_0159_),
    .X(net180));
 sky130_fd_sc_hd__buf_1 fanout181 (.A(_0159_),
    .X(net181));
 sky130_fd_sc_hd__buf_1 fanout182 (.A(net183),
    .X(net182));
 sky130_fd_sc_hd__buf_1 fanout183 (.A(_0156_),
    .X(net183));
 sky130_fd_sc_hd__buf_1 fanout184 (.A(_0154_),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_1 fanout185 (.A(_0154_),
    .X(net185));
 sky130_fd_sc_hd__buf_1 fanout186 (.A(net188),
    .X(net186));
 sky130_fd_sc_hd__clkbuf_1 fanout187 (.A(net188),
    .X(net187));
 sky130_fd_sc_hd__buf_1 fanout188 (.A(_0153_),
    .X(net188));
 sky130_fd_sc_hd__buf_1 fanout189 (.A(net190),
    .X(net189));
 sky130_fd_sc_hd__buf_1 fanout190 (.A(_0152_),
    .X(net190));
 sky130_fd_sc_hd__buf_1 fanout191 (.A(_0146_),
    .X(net191));
 sky130_fd_sc_hd__buf_1 fanout192 (.A(_0146_),
    .X(net192));
 sky130_fd_sc_hd__buf_1 fanout193 (.A(_0145_),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_1 fanout194 (.A(_0145_),
    .X(net194));
 sky130_fd_sc_hd__buf_1 fanout195 (.A(net196),
    .X(net195));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout196 (.A(_0144_),
    .X(net196));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout197 (.A(_0143_),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_1 fanout198 (.A(_0143_),
    .X(net198));
 sky130_fd_sc_hd__buf_1 fanout199 (.A(net200),
    .X(net199));
 sky130_fd_sc_hd__buf_1 fanout200 (.A(net201),
    .X(net200));
 sky130_fd_sc_hd__clkbuf_2 fanout201 (.A(_0141_),
    .X(net201));
 sky130_fd_sc_hd__buf_1 fanout202 (.A(_0140_),
    .X(net202));
 sky130_fd_sc_hd__clkbuf_1 fanout203 (.A(net204),
    .X(net203));
 sky130_fd_sc_hd__clkbuf_2 fanout204 (.A(_0140_),
    .X(net204));
 sky130_fd_sc_hd__buf_1 fanout205 (.A(_0139_),
    .X(net205));
 sky130_fd_sc_hd__buf_1 fanout206 (.A(_0138_),
    .X(net206));
 sky130_fd_sc_hd__clkbuf_1 fanout207 (.A(_0138_),
    .X(net207));
 sky130_fd_sc_hd__buf_1 fanout208 (.A(_0137_),
    .X(net208));
 sky130_fd_sc_hd__buf_1 fanout209 (.A(_0137_),
    .X(net209));
 sky130_fd_sc_hd__buf_1 fanout210 (.A(net211),
    .X(net210));
 sky130_fd_sc_hd__buf_1 fanout211 (.A(_0134_),
    .X(net211));
 sky130_fd_sc_hd__buf_1 fanout212 (.A(_0132_),
    .X(net212));
 sky130_fd_sc_hd__buf_1 fanout213 (.A(net214),
    .X(net213));
 sky130_fd_sc_hd__clkbuf_2 fanout214 (.A(_0132_),
    .X(net214));
 sky130_fd_sc_hd__buf_1 fanout215 (.A(_0131_),
    .X(net215));
 sky130_fd_sc_hd__clkbuf_1 fanout216 (.A(net217),
    .X(net216));
 sky130_fd_sc_hd__clkbuf_2 fanout217 (.A(_0131_),
    .X(net217));
 sky130_fd_sc_hd__buf_1 fanout218 (.A(_0127_),
    .X(net218));
 sky130_fd_sc_hd__clkbuf_1 fanout219 (.A(_0127_),
    .X(net219));
 sky130_fd_sc_hd__buf_1 fanout220 (.A(net222),
    .X(net220));
 sky130_fd_sc_hd__clkbuf_1 fanout221 (.A(net222),
    .X(net221));
 sky130_fd_sc_hd__clkbuf_2 fanout222 (.A(_0126_),
    .X(net222));
 sky130_fd_sc_hd__buf_1 fanout223 (.A(_0125_),
    .X(net223));
 sky130_fd_sc_hd__buf_1 fanout224 (.A(_0125_),
    .X(net224));
 sky130_fd_sc_hd__buf_1 fanout225 (.A(net227),
    .X(net225));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout226 (.A(net227),
    .X(net226));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout227 (.A(_0124_),
    .X(net227));
 sky130_fd_sc_hd__buf_1 fanout228 (.A(net229),
    .X(net228));
 sky130_fd_sc_hd__buf_1 fanout229 (.A(net230),
    .X(net229));
 sky130_fd_sc_hd__clkbuf_2 fanout230 (.A(_0121_),
    .X(net230));
 sky130_fd_sc_hd__buf_1 fanout231 (.A(_0120_),
    .X(net231));
 sky130_fd_sc_hd__buf_1 fanout232 (.A(_0120_),
    .X(net232));
 sky130_fd_sc_hd__buf_1 fanout233 (.A(_0119_),
    .X(net233));
 sky130_fd_sc_hd__buf_1 fanout234 (.A(net235),
    .X(net234));
 sky130_fd_sc_hd__buf_1 fanout235 (.A(_0119_),
    .X(net235));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout236 (.A(_0118_),
    .X(net236));
 sky130_fd_sc_hd__buf_1 fanout237 (.A(_0118_),
    .X(net237));
 sky130_fd_sc_hd__buf_1 fanout238 (.A(net239),
    .X(net238));
 sky130_fd_sc_hd__clkbuf_2 fanout239 (.A(_0111_),
    .X(net239));
 sky130_fd_sc_hd__buf_1 fanout240 (.A(_0109_),
    .X(net240));
 sky130_fd_sc_hd__clkbuf_1 fanout241 (.A(_0109_),
    .X(net241));
 sky130_fd_sc_hd__buf_1 fanout242 (.A(net243),
    .X(net242));
 sky130_fd_sc_hd__buf_1 fanout243 (.A(_0108_),
    .X(net243));
 sky130_fd_sc_hd__buf_1 fanout244 (.A(_0105_),
    .X(net244));
 sky130_fd_sc_hd__clkbuf_1 fanout245 (.A(_0105_),
    .X(net245));
 sky130_fd_sc_hd__buf_1 fanout246 (.A(_0104_),
    .X(net246));
 sky130_fd_sc_hd__buf_1 fanout247 (.A(_0104_),
    .X(net247));
 sky130_fd_sc_hd__buf_1 fanout248 (.A(_0102_),
    .X(net248));
 sky130_fd_sc_hd__clkbuf_1 fanout249 (.A(_0102_),
    .X(net249));
 sky130_fd_sc_hd__buf_1 fanout250 (.A(net251),
    .X(net250));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout251 (.A(_0101_),
    .X(net251));
 sky130_fd_sc_hd__buf_1 fanout252 (.A(_0095_),
    .X(net252));
 sky130_fd_sc_hd__clkbuf_1 fanout253 (.A(_0095_),
    .X(net253));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout254 (.A(_0094_),
    .X(net254));
 sky130_fd_sc_hd__clkbuf_1 fanout255 (.A(_0094_),
    .X(net255));
 sky130_fd_sc_hd__clkbuf_2 fanout256 (.A(_0092_),
    .X(net256));
 sky130_fd_sc_hd__clkbuf_1 fanout257 (.A(_0092_),
    .X(net257));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout258 (.A(_0091_),
    .X(net258));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout259 (.A(_0091_),
    .X(net259));
 sky130_fd_sc_hd__buf_1 fanout260 (.A(net261),
    .X(net260));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout261 (.A(_0087_),
    .X(net261));
 sky130_fd_sc_hd__buf_1 fanout262 (.A(net263),
    .X(net262));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout263 (.A(_0086_),
    .X(net263));
 sky130_fd_sc_hd__buf_1 fanout264 (.A(_0085_),
    .X(net264));
 sky130_fd_sc_hd__clkbuf_1 fanout265 (.A(_0085_),
    .X(net265));
 sky130_fd_sc_hd__buf_1 fanout266 (.A(_0084_),
    .X(net266));
 sky130_fd_sc_hd__buf_1 fanout267 (.A(_0084_),
    .X(net267));
 sky130_fd_sc_hd__buf_1 fanout268 (.A(_0079_),
    .X(net268));
 sky130_fd_sc_hd__clkbuf_1 fanout269 (.A(_0079_),
    .X(net269));
 sky130_fd_sc_hd__buf_1 fanout270 (.A(_0078_),
    .X(net270));
 sky130_fd_sc_hd__buf_1 fanout271 (.A(_0077_),
    .X(net271));
 sky130_fd_sc_hd__buf_1 fanout272 (.A(net274),
    .X(net272));
 sky130_fd_sc_hd__clkbuf_1 fanout273 (.A(net274),
    .X(net273));
 sky130_fd_sc_hd__buf_1 fanout274 (.A(net275),
    .X(net274));
 sky130_fd_sc_hd__buf_1 fanout275 (.A(_0076_),
    .X(net275));
 sky130_fd_sc_hd__buf_1 fanout276 (.A(net277),
    .X(net276));
 sky130_fd_sc_hd__buf_1 fanout277 (.A(_0072_),
    .X(net277));
 sky130_fd_sc_hd__buf_1 fanout278 (.A(_0071_),
    .X(net278));
 sky130_fd_sc_hd__buf_1 fanout279 (.A(_0070_),
    .X(net279));
 sky130_fd_sc_hd__buf_1 fanout280 (.A(net281),
    .X(net280));
 sky130_fd_sc_hd__buf_1 fanout281 (.A(_0069_),
    .X(net281));
 sky130_fd_sc_hd__buf_1 fanout282 (.A(net284),
    .X(net282));
 sky130_fd_sc_hd__clkbuf_1 fanout283 (.A(net284),
    .X(net283));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout284 (.A(_0065_),
    .X(net284));
 sky130_fd_sc_hd__buf_1 fanout285 (.A(net286),
    .X(net285));
 sky130_fd_sc_hd__buf_1 fanout286 (.A(_0063_),
    .X(net286));
 sky130_fd_sc_hd__buf_1 fanout287 (.A(_0062_),
    .X(net287));
 sky130_fd_sc_hd__buf_1 fanout288 (.A(_0057_),
    .X(net288));
 sky130_fd_sc_hd__buf_1 fanout289 (.A(_0057_),
    .X(net289));
 sky130_fd_sc_hd__buf_1 fanout290 (.A(net291),
    .X(net290));
 sky130_fd_sc_hd__clkbuf_2 fanout291 (.A(_0056_),
    .X(net291));
 sky130_fd_sc_hd__buf_1 fanout292 (.A(_0055_),
    .X(net292));
 sky130_fd_sc_hd__buf_1 fanout293 (.A(_0055_),
    .X(net293));
 sky130_fd_sc_hd__buf_1 fanout294 (.A(_0054_),
    .X(net294));
 sky130_fd_sc_hd__clkbuf_1 fanout295 (.A(_0054_),
    .X(net295));
 sky130_fd_sc_hd__buf_1 fanout296 (.A(net297),
    .X(net296));
 sky130_fd_sc_hd__buf_1 fanout297 (.A(net298),
    .X(net297));
 sky130_fd_sc_hd__buf_1 fanout298 (.A(net299),
    .X(net298));
 sky130_fd_sc_hd__buf_1 fanout299 (.A(_0046_),
    .X(net299));
 sky130_fd_sc_hd__buf_1 fanout300 (.A(net302),
    .X(net300));
 sky130_fd_sc_hd__clkbuf_1 fanout301 (.A(net302),
    .X(net301));
 sky130_fd_sc_hd__buf_1 fanout302 (.A(net303),
    .X(net302));
 sky130_fd_sc_hd__buf_1 fanout303 (.A(_0045_),
    .X(net303));
 sky130_fd_sc_hd__buf_1 fanout304 (.A(_0044_),
    .X(net304));
 sky130_fd_sc_hd__buf_1 fanout305 (.A(net306),
    .X(net305));
 sky130_fd_sc_hd__buf_1 fanout306 (.A(_0043_),
    .X(net306));
 sky130_fd_sc_hd__buf_1 fanout307 (.A(net308),
    .X(net307));
 sky130_fd_sc_hd__buf_1 fanout308 (.A(_0039_),
    .X(net308));
 sky130_fd_sc_hd__buf_1 fanout309 (.A(_0038_),
    .X(net309));
 sky130_fd_sc_hd__buf_1 fanout310 (.A(net311),
    .X(net310));
 sky130_fd_sc_hd__buf_1 fanout311 (.A(_0037_),
    .X(net311));
 sky130_fd_sc_hd__buf_1 fanout312 (.A(_0036_),
    .X(net312));
 sky130_fd_sc_hd__clkbuf_2 fanout313 (.A(net314),
    .X(net313));
 sky130_fd_sc_hd__clkbuf_2 fanout314 (.A(_0690_),
    .X(net314));
 sky130_fd_sc_hd__buf_1 fanout315 (.A(_0687_),
    .X(net315));
 sky130_fd_sc_hd__clkbuf_1 fanout316 (.A(net317),
    .X(net316));
 sky130_fd_sc_hd__buf_1 max_cap317 (.A(_0687_),
    .X(net317));
 sky130_fd_sc_hd__buf_1 fanout318 (.A(net319),
    .X(net318));
 sky130_fd_sc_hd__clkbuf_1 fanout319 (.A(net320),
    .X(net319));
 sky130_fd_sc_hd__clkbuf_1 fanout320 (.A(net321),
    .X(net320));
 sky130_fd_sc_hd__buf_1 fanout321 (.A(_0684_),
    .X(net321));
 sky130_fd_sc_hd__buf_1 fanout322 (.A(_0681_),
    .X(net322));
 sky130_fd_sc_hd__clkbuf_1 fanout323 (.A(_0681_),
    .X(net323));
 sky130_fd_sc_hd__buf_1 fanout324 (.A(_0676_),
    .X(net324));
 sky130_fd_sc_hd__clkbuf_1 fanout325 (.A(net326),
    .X(net325));
 sky130_fd_sc_hd__clkbuf_2 fanout326 (.A(_0676_),
    .X(net326));
 sky130_fd_sc_hd__buf_1 fanout327 (.A(net329),
    .X(net327));
 sky130_fd_sc_hd__clkbuf_1 fanout328 (.A(net329),
    .X(net328));
 sky130_fd_sc_hd__clkbuf_1 fanout329 (.A(net330),
    .X(net329));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout330 (.A(_0674_),
    .X(net330));
 sky130_fd_sc_hd__clkbuf_2 fanout331 (.A(_0671_),
    .X(net331));
 sky130_fd_sc_hd__clkbuf_1 fanout332 (.A(_0671_),
    .X(net332));
 sky130_fd_sc_hd__clkbuf_2 fanout333 (.A(_0668_),
    .X(net333));
 sky130_fd_sc_hd__buf_1 fanout334 (.A(_0668_),
    .X(net334));
 sky130_fd_sc_hd__buf_1 fanout335 (.A(net337),
    .X(net335));
 sky130_fd_sc_hd__clkbuf_1 fanout336 (.A(net337),
    .X(net336));
 sky130_fd_sc_hd__buf_1 fanout337 (.A(net341),
    .X(net337));
 sky130_fd_sc_hd__buf_1 fanout338 (.A(net340),
    .X(net338));
 sky130_fd_sc_hd__buf_1 fanout339 (.A(net340),
    .X(net339));
 sky130_fd_sc_hd__buf_1 fanout340 (.A(net341),
    .X(net340));
 sky130_fd_sc_hd__buf_1 fanout341 (.A(_0184_),
    .X(net341));
 sky130_fd_sc_hd__buf_1 fanout342 (.A(net343),
    .X(net342));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout343 (.A(net347),
    .X(net343));
 sky130_fd_sc_hd__buf_1 fanout344 (.A(net345),
    .X(net344));
 sky130_fd_sc_hd__buf_1 fanout345 (.A(net346),
    .X(net345));
 sky130_fd_sc_hd__buf_1 fanout346 (.A(net347),
    .X(net346));
 sky130_fd_sc_hd__buf_1 fanout347 (.A(_0177_),
    .X(net347));
 sky130_fd_sc_hd__buf_1 fanout348 (.A(net349),
    .X(net348));
 sky130_fd_sc_hd__buf_1 fanout349 (.A(net353),
    .X(net349));
 sky130_fd_sc_hd__buf_1 fanout350 (.A(net351),
    .X(net350));
 sky130_fd_sc_hd__buf_1 fanout351 (.A(net352),
    .X(net351));
 sky130_fd_sc_hd__clkbuf_1 fanout352 (.A(net353),
    .X(net352));
 sky130_fd_sc_hd__buf_1 fanout353 (.A(net354),
    .X(net353));
 sky130_fd_sc_hd__buf_1 fanout354 (.A(_0151_),
    .X(net354));
 sky130_fd_sc_hd__buf_1 fanout355 (.A(net359),
    .X(net355));
 sky130_fd_sc_hd__buf_1 fanout356 (.A(net357),
    .X(net356));
 sky130_fd_sc_hd__buf_1 fanout357 (.A(net358),
    .X(net357));
 sky130_fd_sc_hd__clkbuf_1 fanout358 (.A(net359),
    .X(net358));
 sky130_fd_sc_hd__buf_1 fanout359 (.A(net360),
    .X(net359));
 sky130_fd_sc_hd__buf_1 fanout360 (.A(_0150_),
    .X(net360));
 sky130_fd_sc_hd__buf_1 fanout361 (.A(net366),
    .X(net361));
 sky130_fd_sc_hd__buf_1 fanout362 (.A(net366),
    .X(net362));
 sky130_fd_sc_hd__buf_1 fanout363 (.A(net366),
    .X(net363));
 sky130_fd_sc_hd__clkbuf_1 fanout364 (.A(net365),
    .X(net364));
 sky130_fd_sc_hd__buf_1 fanout365 (.A(net366),
    .X(net365));
 sky130_fd_sc_hd__buf_1 fanout366 (.A(_0117_),
    .X(net366));
 sky130_fd_sc_hd__buf_1 fanout367 (.A(net372),
    .X(net367));
 sky130_fd_sc_hd__buf_1 fanout368 (.A(net372),
    .X(net368));
 sky130_fd_sc_hd__buf_1 fanout369 (.A(net372),
    .X(net369));
 sky130_fd_sc_hd__clkbuf_1 fanout370 (.A(net371),
    .X(net370));
 sky130_fd_sc_hd__buf_1 fanout371 (.A(net372),
    .X(net371));
 sky130_fd_sc_hd__buf_1 fanout372 (.A(_0116_),
    .X(net372));
 sky130_fd_sc_hd__buf_1 fanout373 (.A(net374),
    .X(net373));
 sky130_fd_sc_hd__buf_1 fanout374 (.A(net375),
    .X(net374));
 sky130_fd_sc_hd__buf_1 fanout375 (.A(net376),
    .X(net375));
 sky130_fd_sc_hd__buf_1 fanout376 (.A(net378),
    .X(net376));
 sky130_fd_sc_hd__buf_1 fanout377 (.A(_0100_),
    .X(net377));
 sky130_fd_sc_hd__clkbuf_1 fanout378 (.A(_0100_),
    .X(net378));
 sky130_fd_sc_hd__buf_1 fanout379 (.A(net380),
    .X(net379));
 sky130_fd_sc_hd__buf_1 fanout380 (.A(net381),
    .X(net380));
 sky130_fd_sc_hd__buf_1 fanout381 (.A(net382),
    .X(net381));
 sky130_fd_sc_hd__buf_1 fanout382 (.A(net383),
    .X(net382));
 sky130_fd_sc_hd__buf_1 fanout383 (.A(net385),
    .X(net383));
 sky130_fd_sc_hd__clkbuf_1 wire384 (.A(_0099_),
    .X(net384));
 sky130_fd_sc_hd__clkbuf_1 max_cap385 (.A(_0099_),
    .X(net385));
 sky130_fd_sc_hd__buf_1 fanout386 (.A(net391),
    .X(net386));
 sky130_fd_sc_hd__buf_1 fanout387 (.A(net388),
    .X(net387));
 sky130_fd_sc_hd__buf_1 fanout388 (.A(net389),
    .X(net388));
 sky130_fd_sc_hd__clkbuf_1 fanout389 (.A(net390),
    .X(net389));
 sky130_fd_sc_hd__buf_1 fanout390 (.A(net391),
    .X(net390));
 sky130_fd_sc_hd__buf_1 fanout391 (.A(_0083_),
    .X(net391));
 sky130_fd_sc_hd__buf_1 fanout392 (.A(net397),
    .X(net392));
 sky130_fd_sc_hd__buf_1 fanout393 (.A(net394),
    .X(net393));
 sky130_fd_sc_hd__buf_1 fanout394 (.A(net395),
    .X(net394));
 sky130_fd_sc_hd__clkbuf_1 fanout395 (.A(net396),
    .X(net395));
 sky130_fd_sc_hd__buf_1 fanout396 (.A(net397),
    .X(net396));
 sky130_fd_sc_hd__buf_1 fanout397 (.A(_0082_),
    .X(net397));
 sky130_fd_sc_hd__buf_1 fanout398 (.A(net399),
    .X(net398));
 sky130_fd_sc_hd__buf_1 fanout399 (.A(net405),
    .X(net399));
 sky130_fd_sc_hd__buf_1 fanout400 (.A(net401),
    .X(net400));
 sky130_fd_sc_hd__clkbuf_1 fanout401 (.A(net402),
    .X(net401));
 sky130_fd_sc_hd__buf_1 fanout402 (.A(net403),
    .X(net402));
 sky130_fd_sc_hd__buf_1 fanout403 (.A(net404),
    .X(net403));
 sky130_fd_sc_hd__buf_1 fanout404 (.A(net405),
    .X(net404));
 sky130_fd_sc_hd__clkbuf_1 fanout405 (.A(_0068_),
    .X(net405));
 sky130_fd_sc_hd__buf_1 fanout406 (.A(net408),
    .X(net406));
 sky130_fd_sc_hd__clkbuf_1 fanout407 (.A(net408),
    .X(net407));
 sky130_fd_sc_hd__buf_1 fanout408 (.A(net414),
    .X(net408));
 sky130_fd_sc_hd__buf_1 fanout409 (.A(net410),
    .X(net409));
 sky130_fd_sc_hd__buf_1 fanout410 (.A(net411),
    .X(net410));
 sky130_fd_sc_hd__clkbuf_1 fanout411 (.A(net412),
    .X(net411));
 sky130_fd_sc_hd__clkbuf_1 fanout412 (.A(net413),
    .X(net412));
 sky130_fd_sc_hd__buf_1 fanout413 (.A(net414),
    .X(net413));
 sky130_fd_sc_hd__clkbuf_1 fanout414 (.A(_0067_),
    .X(net414));
 sky130_fd_sc_hd__buf_1 fanout415 (.A(net416),
    .X(net415));
 sky130_fd_sc_hd__buf_1 fanout416 (.A(net417),
    .X(net416));
 sky130_fd_sc_hd__clkbuf_1 fanout417 (.A(net418),
    .X(net417));
 sky130_fd_sc_hd__buf_1 fanout418 (.A(net421),
    .X(net418));
 sky130_fd_sc_hd__buf_1 fanout419 (.A(net420),
    .X(net419));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout420 (.A(net421),
    .X(net420));
 sky130_fd_sc_hd__buf_1 fanout421 (.A(_0053_),
    .X(net421));
 sky130_fd_sc_hd__buf_1 fanout422 (.A(net423),
    .X(net422));
 sky130_fd_sc_hd__buf_1 fanout423 (.A(net424),
    .X(net423));
 sky130_fd_sc_hd__clkbuf_1 fanout424 (.A(net425),
    .X(net424));
 sky130_fd_sc_hd__buf_1 fanout425 (.A(net428),
    .X(net425));
 sky130_fd_sc_hd__buf_1 fanout426 (.A(net428),
    .X(net426));
 sky130_fd_sc_hd__buf_1 fanout427 (.A(net428),
    .X(net427));
 sky130_fd_sc_hd__buf_1 fanout428 (.A(_0052_),
    .X(net428));
 sky130_fd_sc_hd__buf_1 fanout429 (.A(net431),
    .X(net429));
 sky130_fd_sc_hd__clkbuf_1 fanout430 (.A(net431),
    .X(net430));
 sky130_fd_sc_hd__buf_1 fanout431 (.A(net435),
    .X(net431));
 sky130_fd_sc_hd__buf_1 fanout432 (.A(net433),
    .X(net432));
 sky130_fd_sc_hd__buf_1 fanout433 (.A(net434),
    .X(net433));
 sky130_fd_sc_hd__buf_1 fanout434 (.A(net435),
    .X(net434));
 sky130_fd_sc_hd__buf_1 fanout435 (.A(_0035_),
    .X(net435));
 sky130_fd_sc_hd__buf_1 fanout436 (.A(net438),
    .X(net436));
 sky130_fd_sc_hd__clkbuf_1 fanout437 (.A(net438),
    .X(net437));
 sky130_fd_sc_hd__buf_1 fanout438 (.A(net442),
    .X(net438));
 sky130_fd_sc_hd__buf_1 fanout439 (.A(net440),
    .X(net439));
 sky130_fd_sc_hd__buf_1 fanout440 (.A(net441),
    .X(net440));
 sky130_fd_sc_hd__buf_1 fanout441 (.A(net442),
    .X(net441));
 sky130_fd_sc_hd__buf_1 fanout442 (.A(_0034_),
    .X(net442));
 sky130_fd_sc_hd__buf_1 fanout443 (.A(net445),
    .X(net443));
 sky130_fd_sc_hd__buf_1 fanout444 (.A(net445),
    .X(net444));
 sky130_fd_sc_hd__clkbuf_1 fanout445 (.A(net446),
    .X(net445));
 sky130_fd_sc_hd__buf_1 fanout446 (.A(net449),
    .X(net446));
 sky130_fd_sc_hd__buf_1 fanout447 (.A(net448),
    .X(net447));
 sky130_fd_sc_hd__buf_1 fanout448 (.A(net449),
    .X(net448));
 sky130_fd_sc_hd__buf_1 fanout449 (.A(_0689_),
    .X(net449));
 sky130_fd_sc_hd__buf_1 fanout450 (.A(net452),
    .X(net450));
 sky130_fd_sc_hd__buf_1 fanout451 (.A(net452),
    .X(net451));
 sky130_fd_sc_hd__clkbuf_1 fanout452 (.A(net453),
    .X(net452));
 sky130_fd_sc_hd__buf_1 fanout453 (.A(net456),
    .X(net453));
 sky130_fd_sc_hd__buf_1 fanout454 (.A(net455),
    .X(net454));
 sky130_fd_sc_hd__buf_1 fanout455 (.A(net456),
    .X(net455));
 sky130_fd_sc_hd__buf_1 fanout456 (.A(_0688_),
    .X(net456));
 sky130_fd_sc_hd__buf_1 fanout457 (.A(_0686_),
    .X(net457));
 sky130_fd_sc_hd__buf_1 fanout458 (.A(_0686_),
    .X(net458));
 sky130_fd_sc_hd__buf_1 fanout459 (.A(net460),
    .X(net459));
 sky130_fd_sc_hd__buf_1 fanout460 (.A(net461),
    .X(net460));
 sky130_fd_sc_hd__buf_1 fanout461 (.A(net466),
    .X(net461));
 sky130_fd_sc_hd__buf_1 fanout462 (.A(net463),
    .X(net462));
 sky130_fd_sc_hd__clkbuf_1 fanout463 (.A(net464),
    .X(net463));
 sky130_fd_sc_hd__buf_1 fanout464 (.A(net465),
    .X(net464));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout465 (.A(net466),
    .X(net465));
 sky130_fd_sc_hd__buf_1 fanout466 (.A(_0683_),
    .X(net466));
 sky130_fd_sc_hd__buf_1 fanout467 (.A(net468),
    .X(net467));
 sky130_fd_sc_hd__buf_1 fanout468 (.A(net469),
    .X(net468));
 sky130_fd_sc_hd__buf_1 fanout469 (.A(net474),
    .X(net469));
 sky130_fd_sc_hd__buf_1 fanout470 (.A(net471),
    .X(net470));
 sky130_fd_sc_hd__clkbuf_1 fanout471 (.A(net472),
    .X(net471));
 sky130_fd_sc_hd__buf_1 fanout472 (.A(net473),
    .X(net472));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout473 (.A(net474),
    .X(net473));
 sky130_fd_sc_hd__buf_1 fanout474 (.A(_0682_),
    .X(net474));
 sky130_fd_sc_hd__buf_1 fanout475 (.A(net476),
    .X(net475));
 sky130_fd_sc_hd__buf_1 fanout476 (.A(net477),
    .X(net476));
 sky130_fd_sc_hd__buf_1 fanout477 (.A(net481),
    .X(net477));
 sky130_fd_sc_hd__buf_1 fanout478 (.A(net480),
    .X(net478));
 sky130_fd_sc_hd__clkbuf_1 fanout479 (.A(net480),
    .X(net479));
 sky130_fd_sc_hd__clkbuf_1 fanout480 (.A(net481),
    .X(net480));
 sky130_fd_sc_hd__buf_1 fanout481 (.A(_0680_),
    .X(net481));
 sky130_fd_sc_hd__buf_1 fanout482 (.A(net483),
    .X(net482));
 sky130_fd_sc_hd__buf_1 fanout483 (.A(net484),
    .X(net483));
 sky130_fd_sc_hd__buf_1 fanout484 (.A(net488),
    .X(net484));
 sky130_fd_sc_hd__buf_1 fanout485 (.A(net487),
    .X(net485));
 sky130_fd_sc_hd__clkbuf_1 fanout486 (.A(net487),
    .X(net486));
 sky130_fd_sc_hd__clkbuf_1 fanout487 (.A(net488),
    .X(net487));
 sky130_fd_sc_hd__buf_1 fanout488 (.A(_0679_),
    .X(net488));
 sky130_fd_sc_hd__buf_1 fanout489 (.A(_0675_),
    .X(net489));
 sky130_fd_sc_hd__buf_1 fanout490 (.A(_0675_),
    .X(net490));
 sky130_fd_sc_hd__buf_1 fanout491 (.A(net492),
    .X(net491));
 sky130_fd_sc_hd__buf_1 fanout492 (.A(net493),
    .X(net492));
 sky130_fd_sc_hd__clkbuf_1 fanout493 (.A(net494),
    .X(net493));
 sky130_fd_sc_hd__clkbuf_1 fanout494 (.A(net496),
    .X(net494));
 sky130_fd_sc_hd__buf_1 fanout495 (.A(net496),
    .X(net495));
 sky130_fd_sc_hd__buf_1 fanout496 (.A(_0673_),
    .X(net496));
 sky130_fd_sc_hd__clkbuf_1 fanout497 (.A(_0673_),
    .X(net497));
 sky130_fd_sc_hd__buf_1 fanout498 (.A(net502),
    .X(net498));
 sky130_fd_sc_hd__buf_1 fanout499 (.A(net500),
    .X(net499));
 sky130_fd_sc_hd__buf_1 fanout500 (.A(net501),
    .X(net500));
 sky130_fd_sc_hd__clkbuf_1 fanout501 (.A(net502),
    .X(net501));
 sky130_fd_sc_hd__buf_1 fanout502 (.A(net503),
    .X(net502));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout503 (.A(_0672_),
    .X(net503));
 sky130_fd_sc_hd__buf_1 fanout504 (.A(net505),
    .X(net504));
 sky130_fd_sc_hd__buf_1 fanout505 (.A(net506),
    .X(net505));
 sky130_fd_sc_hd__clkbuf_1 fanout506 (.A(net507),
    .X(net506));
 sky130_fd_sc_hd__buf_1 fanout507 (.A(net510),
    .X(net507));
 sky130_fd_sc_hd__buf_1 fanout508 (.A(net509),
    .X(net508));
 sky130_fd_sc_hd__buf_1 fanout509 (.A(net510),
    .X(net509));
 sky130_fd_sc_hd__buf_1 fanout510 (.A(_0670_),
    .X(net510));
 sky130_fd_sc_hd__buf_1 fanout511 (.A(net512),
    .X(net511));
 sky130_fd_sc_hd__buf_1 fanout512 (.A(net513),
    .X(net512));
 sky130_fd_sc_hd__clkbuf_1 fanout513 (.A(net514),
    .X(net513));
 sky130_fd_sc_hd__buf_1 fanout514 (.A(net517),
    .X(net514));
 sky130_fd_sc_hd__buf_1 fanout515 (.A(net516),
    .X(net515));
 sky130_fd_sc_hd__buf_1 fanout516 (.A(net517),
    .X(net516));
 sky130_fd_sc_hd__buf_1 fanout517 (.A(_0669_),
    .X(net517));
 sky130_fd_sc_hd__buf_1 fanout518 (.A(net522),
    .X(net518));
 sky130_fd_sc_hd__buf_1 fanout519 (.A(net522),
    .X(net519));
 sky130_fd_sc_hd__buf_1 fanout520 (.A(net522),
    .X(net520));
 sky130_fd_sc_hd__buf_1 fanout521 (.A(net522),
    .X(net521));
 sky130_fd_sc_hd__buf_1 fanout522 (.A(_0666_),
    .X(net522));
 sky130_fd_sc_hd__buf_1 fanout523 (.A(net524),
    .X(net523));
 sky130_fd_sc_hd__buf_1 fanout524 (.A(net525),
    .X(net524));
 sky130_fd_sc_hd__clkbuf_1 fanout525 (.A(net526),
    .X(net525));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout526 (.A(net529),
    .X(net526));
 sky130_fd_sc_hd__buf_1 fanout527 (.A(net529),
    .X(net527));
 sky130_fd_sc_hd__clkbuf_1 fanout528 (.A(net529),
    .X(net528));
 sky130_fd_sc_hd__buf_1 fanout529 (.A(_0658_),
    .X(net529));
 sky130_fd_sc_hd__buf_1 fanout530 (.A(net531),
    .X(net530));
 sky130_fd_sc_hd__buf_1 fanout531 (.A(net534),
    .X(net531));
 sky130_fd_sc_hd__buf_1 fanout532 (.A(net534),
    .X(net532));
 sky130_fd_sc_hd__buf_1 fanout533 (.A(net534),
    .X(net533));
 sky130_fd_sc_hd__buf_1 fanout534 (.A(_0648_),
    .X(net534));
 sky130_fd_sc_hd__buf_1 fanout535 (.A(net536),
    .X(net535));
 sky130_fd_sc_hd__buf_1 fanout536 (.A(net537),
    .X(net536));
 sky130_fd_sc_hd__clkbuf_1 fanout537 (.A(net538),
    .X(net537));
 sky130_fd_sc_hd__buf_1 fanout538 (.A(net541),
    .X(net538));
 sky130_fd_sc_hd__buf_1 fanout539 (.A(net541),
    .X(net539));
 sky130_fd_sc_hd__clkbuf_1 fanout540 (.A(net541),
    .X(net540));
 sky130_fd_sc_hd__buf_1 fanout541 (.A(_0638_),
    .X(net541));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout542 (.A(net546),
    .X(net542));
 sky130_fd_sc_hd__buf_1 fanout543 (.A(net545),
    .X(net543));
 sky130_fd_sc_hd__clkbuf_1 fanout544 (.A(net545),
    .X(net544));
 sky130_fd_sc_hd__clkbuf_1 fanout545 (.A(net546),
    .X(net545));
 sky130_fd_sc_hd__buf_1 fanout546 (.A(net547),
    .X(net546));
 sky130_fd_sc_hd__clkbuf_2 fanout547 (.A(net557),
    .X(net547));
 sky130_fd_sc_hd__buf_1 fanout548 (.A(net549),
    .X(net548));
 sky130_fd_sc_hd__clkbuf_1 fanout549 (.A(net556),
    .X(net549));
 sky130_fd_sc_hd__buf_1 fanout550 (.A(net552),
    .X(net550));
 sky130_fd_sc_hd__clkbuf_1 fanout551 (.A(net552),
    .X(net551));
 sky130_fd_sc_hd__clkbuf_1 fanout552 (.A(net555),
    .X(net552));
 sky130_fd_sc_hd__buf_1 fanout553 (.A(net554),
    .X(net553));
 sky130_fd_sc_hd__buf_1 fanout554 (.A(net555),
    .X(net554));
 sky130_fd_sc_hd__buf_1 fanout555 (.A(net556),
    .X(net555));
 sky130_fd_sc_hd__clkbuf_1 fanout556 (.A(net557),
    .X(net556));
 sky130_fd_sc_hd__buf_1 fanout557 (.A(_0628_),
    .X(net557));
 sky130_fd_sc_hd__buf_1 fanout558 (.A(net559),
    .X(net558));
 sky130_fd_sc_hd__clkbuf_1 fanout559 (.A(net563),
    .X(net559));
 sky130_fd_sc_hd__buf_1 fanout560 (.A(net563),
    .X(net560));
 sky130_fd_sc_hd__buf_1 fanout561 (.A(net563),
    .X(net561));
 sky130_fd_sc_hd__clkbuf_1 fanout562 (.A(net563),
    .X(net562));
 sky130_fd_sc_hd__buf_1 fanout563 (.A(\addr0_reg[7] ),
    .X(net563));
 sky130_fd_sc_hd__clkbuf_1 fanout564 (.A(net565),
    .X(net564));
 sky130_fd_sc_hd__clkbuf_1 fanout565 (.A(net569),
    .X(net565));
 sky130_fd_sc_hd__buf_1 fanout566 (.A(net569),
    .X(net566));
 sky130_fd_sc_hd__buf_1 fanout567 (.A(net569),
    .X(net567));
 sky130_fd_sc_hd__clkbuf_1 fanout568 (.A(net569),
    .X(net568));
 sky130_fd_sc_hd__buf_1 fanout569 (.A(\addr0_reg[6] ),
    .X(net569));
 sky130_fd_sc_hd__buf_1 fanout570 (.A(net571),
    .X(net570));
 sky130_fd_sc_hd__clkbuf_1 fanout571 (.A(net572),
    .X(net571));
 sky130_fd_sc_hd__clkbuf_1 fanout572 (.A(net576),
    .X(net572));
 sky130_fd_sc_hd__buf_1 fanout573 (.A(net576),
    .X(net573));
 sky130_fd_sc_hd__buf_1 fanout574 (.A(net575),
    .X(net574));
 sky130_fd_sc_hd__buf_1 fanout575 (.A(net576),
    .X(net575));
 sky130_fd_sc_hd__buf_1 fanout576 (.A(\addr0_reg[5] ),
    .X(net576));
 sky130_fd_sc_hd__buf_1 fanout577 (.A(net578),
    .X(net577));
 sky130_fd_sc_hd__clkbuf_1 fanout578 (.A(net579),
    .X(net578));
 sky130_fd_sc_hd__clkbuf_1 fanout579 (.A(net583),
    .X(net579));
 sky130_fd_sc_hd__buf_1 fanout580 (.A(net583),
    .X(net580));
 sky130_fd_sc_hd__buf_1 fanout581 (.A(net583),
    .X(net581));
 sky130_fd_sc_hd__buf_1 fanout582 (.A(net583),
    .X(net582));
 sky130_fd_sc_hd__buf_1 fanout583 (.A(\addr0_reg[4] ),
    .X(net583));
 sky130_fd_sc_hd__clkbuf_1 fanout584 (.A(net586),
    .X(net584));
 sky130_fd_sc_hd__clkbuf_1 fanout585 (.A(net586),
    .X(net585));
 sky130_fd_sc_hd__clkbuf_1 fanout586 (.A(net587),
    .X(net586));
 sky130_fd_sc_hd__clkbuf_1 fanout587 (.A(net588),
    .X(net587));
 sky130_fd_sc_hd__clkbuf_1 fanout588 (.A(net592),
    .X(net588));
 sky130_fd_sc_hd__buf_1 fanout589 (.A(net590),
    .X(net589));
 sky130_fd_sc_hd__clkbuf_1 fanout590 (.A(net591),
    .X(net590));
 sky130_fd_sc_hd__buf_1 fanout591 (.A(net592),
    .X(net591));
 sky130_fd_sc_hd__clkbuf_1 fanout592 (.A(\addr0_reg[3] ),
    .X(net592));
 sky130_fd_sc_hd__clkbuf_1 fanout593 (.A(net594),
    .X(net593));
 sky130_fd_sc_hd__clkbuf_1 fanout594 (.A(net595),
    .X(net594));
 sky130_fd_sc_hd__clkbuf_1 fanout595 (.A(net596),
    .X(net595));
 sky130_fd_sc_hd__clkbuf_1 fanout596 (.A(net599),
    .X(net596));
 sky130_fd_sc_hd__buf_1 fanout597 (.A(net598),
    .X(net597));
 sky130_fd_sc_hd__buf_1 fanout598 (.A(net599),
    .X(net598));
 sky130_fd_sc_hd__buf_1 fanout599 (.A(\addr0_reg[2] ),
    .X(net599));
 sky130_fd_sc_hd__clkbuf_1 fanout600 (.A(net602),
    .X(net600));
 sky130_fd_sc_hd__clkbuf_1 fanout601 (.A(net602),
    .X(net601));
 sky130_fd_sc_hd__clkbuf_1 fanout602 (.A(net606),
    .X(net602));
 sky130_fd_sc_hd__buf_1 fanout603 (.A(net604),
    .X(net603));
 sky130_fd_sc_hd__clkbuf_1 fanout604 (.A(net605),
    .X(net604));
 sky130_fd_sc_hd__buf_1 fanout605 (.A(net606),
    .X(net605));
 sky130_fd_sc_hd__clkbuf_1 fanout606 (.A(\addr0_reg[1] ),
    .X(net606));
 sky130_fd_sc_hd__clkbuf_1 fanout607 (.A(net609),
    .X(net607));
 sky130_fd_sc_hd__clkbuf_1 fanout608 (.A(net609),
    .X(net608));
 sky130_fd_sc_hd__clkbuf_1 fanout609 (.A(net610),
    .X(net609));
 sky130_fd_sc_hd__clkbuf_1 fanout610 (.A(net611),
    .X(net610));
 sky130_fd_sc_hd__clkbuf_1 fanout611 (.A(net615),
    .X(net611));
 sky130_fd_sc_hd__buf_1 fanout612 (.A(net613),
    .X(net612));
 sky130_fd_sc_hd__clkbuf_1 fanout613 (.A(net614),
    .X(net613));
 sky130_fd_sc_hd__buf_1 fanout614 (.A(net615),
    .X(net614));
 sky130_fd_sc_hd__clkbuf_1 fanout615 (.A(\addr0_reg[0] ),
    .X(net615));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk0 (.A(clk0),
    .X(clknet_0_clk0));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk0 (.A(clknet_0_clk0),
    .X(clknet_2_0__leaf_clk0));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk0 (.A(clknet_0_clk0),
    .X(clknet_2_1__leaf_clk0));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk0 (.A(clknet_0_clk0),
    .X(clknet_2_2__leaf_clk0));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk0 (.A(clknet_0_clk0),
    .X(clknet_2_3__leaf_clk0));
 sky130_fd_sc_hd__bufinv_16 clkload0 (.A(clknet_2_0__leaf_clk0));
 sky130_fd_sc_hd__bufinv_16 clkload1 (.A(clknet_2_1__leaf_clk0));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(net38),
    .X(net616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(net26),
    .X(net617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(net20),
    .X(net618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(net37),
    .X(net619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(net29),
    .X(net620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(net15),
    .X(net621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(net14),
    .X(net622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(net31),
    .X(net623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(net35),
    .X(net624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(net30),
    .X(net625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(net40),
    .X(net626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(net39),
    .X(net627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(net32),
    .X(net628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(net10),
    .X(net629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(net21),
    .X(net630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(net12),
    .X(net631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(net16),
    .X(net632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(net27),
    .X(net633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(net25),
    .X(net634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(net28),
    .X(net635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(net19),
    .X(net636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(net13),
    .X(net637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(net17),
    .X(net638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(net22),
    .X(net639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(net11),
    .X(net640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(net34),
    .X(net641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(net24),
    .X(net642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(net23),
    .X(net643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(net41),
    .X(net644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(net36),
    .X(net645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(net18),
    .X(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_0056_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_0057_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_0060_));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_0105_));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_0123_));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_0140_));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(_0160_));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(_0181_));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_0186_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(_0189_));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(_0192_));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(_0201_));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(_0201_));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(_0201_));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(_0212_));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(_0220_));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(_0220_));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(_0228_));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(_0242_));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(_0249_));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(_0249_));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(_0252_));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(_0281_));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(_0281_));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(_0329_));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(_0344_));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(_0481_));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(_0506_));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(_0527_));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(_0676_));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(clknet_2_1__leaf_clk0));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(_0060_));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(_0094_));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(_0108_));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(_0142_));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(_0255_));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(_0504_));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(_0467_));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(net109));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_18 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_79 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_339 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_6 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_140 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_64 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_22 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_142 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_30 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_143 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_56 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_142 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_341 ();
endmodule
